netcdf no2_conc_rotterdam_20110418_new {
dimensions:
	x = 30 ;
	y = 30 ;
	z = 1 ;
	time = 24 ;
	receptor = 9 ;
	realisation = 7 ;
	dimcrs = 1 ;
variables:
	double x(x) ;
		x:units = "meter" ;
		x:axis = "x" ;
		x:long_name = "x" ;
		x:standard_name = "projection_x_coordinate" ;
	double y(y) ;
		y:units = "meter" ;
		y:axis = "y" ;
		y:long_name = "y" ;
		y:standard_name = "projection_y_coordinate" ;
	double z(z) ;
		z:units = "meter" ;
		z:axis = "z" ;
		z:long_name = "z" ;
		z:standard_name = "height" ;
		z:positive = "up" ;
	int time(time) ;
		time:units = "hours since 2011-04-18 00:00:00 00:00" ;
		time:axis = "t" ;
		time:calendar = "gregorian" ;
		time:long_name = "time" ;
		time:standard_name = "time" ;
	float no2_conc_grid_ctl(time, z, y, x) ;
		no2_conc_grid_ctl:units = "ug m-3" ;
		no2_conc_grid_ctl:missing_value = -9900.f ;
		no2_conc_grid_ctl:long_name = "NO2 main grid concentrations (control)" ;
		no2_conc_grid_ctl:comment = "No comments" ;
		no2_conc_grid_ctl:coordinates = "lat lon" ;
		no2_conc_grid_ctl:_FillValue = -9900.f ;
		no2_conc_grid_ctl:grid_mapping = "crs" ;
		no2_conc_grid_ctl:valid_min = 0.f ;
	int receptor(receptor) ;
		receptor:units = "count" ;
		receptor:long_name = "Receptor indices" ;
	float no2_conc_recp_ctl(time, z, receptor) ;
		no2_conc_recp_ctl:units = "ug m-3" ;
		no2_conc_recp_ctl:missing_value = -9900.f ;
		no2_conc_recp_ctl:long_name = "NO2 receptor concentrations (control)" ;
		no2_conc_recp_ctl:comment = "No comments" ;
		no2_conc_recp_ctl:coordinates = "rlat rlon" ;
		no2_conc_recp_ctl:_FillValue = -9900.f ;
		no2_conc_recp_ctl:valid_min = 0.f ;
	int realisation(realisation) ;
		realisation:units = "count" ;
		realisation:long_name = "realization" ;
		realisation:standard_name = "realization" ;
		realisation:ref = "http://www.uncertml.org/samples/continuous-realisation" ;
	float no2_conc_grid_ens(realisation, time, z, y, x) ;
		no2_conc_grid_ens:units = "ug m-3" ;
		no2_conc_grid_ens:missing_value = -9900.f ;
		no2_conc_grid_ens:long_name = "NO2 main grid concentrations (ensemble)" ;
		no2_conc_grid_ens:comment = "No comments" ;
		no2_conc_grid_ens:coordinates = "lat lon" ;
		no2_conc_grid_ens:_FillValue = -9900.f ;
		no2_conc_grid_ens:grid_mapping = "crs" ;
		no2_conc_grid_ens:valid_min = 0.f ;
		no2_conc_grid_ens:ref = "http://www.uncertml.org/samples/random" ;
	float no2_conc_recp_ens(realisation, time, z, receptor) ;
		no2_conc_recp_ens:units = "ug m-3" ;
		no2_conc_recp_ens:missing_value = -9900.f ;
		no2_conc_recp_ens:long_name = "NO2 receptor concentrations (ensemble)" ;
		no2_conc_recp_ens:comment = "No comments" ;
		no2_conc_recp_ens:coordinates = "rlat rlon" ;
		no2_conc_recp_ens:_FillValue = -9900.f ;
		no2_conc_recp_ens:valid_min = 0.f ;
		no2_conc_recp_ens:ref = "http://www.uncertml.org/samples/random" ;
	int dimcrs(dimcrs) ;
		dimcrs:units = "count" ;
		dimcrs:long_name = "CRS dummy dimension" ;
	char crs(dimcrs) ;
		crs:units = "m" ;
		crs:missing_value = "NA" ;
		crs:_CoordinateTransformType = "Projection" ;
		crs:grid_mapping_name = "transverse_mercator" ;
		crs:proj4string = "+proj=tmerc +lat_0=51.91667 +lon_0=4.475 +k=0.9996 +ellps=WGS84 +units=m" ;
	double lat(y, x) ;
		lat:units = "degrees_north" ;
		lat:missing_value = -9900. ;
		lat:long_name = "Main grid latitudes" ;
		lat:standard_name = "latitude" ;
		lat:valid_min = -90. ;
		lat:valid_max = 90. ;
	double lon(y, x) ;
		lon:units = "degrees_east" ;
		lon:missing_value = -9900. ;
		lon:long_name = "Main grid longitudes" ;
		lon:standard_name = "longitude" ;
		lon:valid_min = -180. ;
		lon:valid_max = 180. ;
	double rlat(receptor) ;
		rlat:units = "degrees_north" ;
		rlat:missing_value = -9900. ;
		rlat:long_name = "Receptor latitudes" ;
		rlat:standard_name = "latitude" ;
		rlat:valid_min = -90. ;
		rlat:valid_max = 90. ;
	double rlon(receptor) ;
		rlon:units = "degrees_east" ;
		rlon:missing_value = -9900. ;
		rlon:long_name = "Receptor longitudes" ;
		rlon:standard_name = "longitude" ;
		rlon:valid_min = -180. ;
		rlon:valid_max = 180. ;
	double weights(realisation) ;
		weights:units = "" ;
		weights:missing_value = -9900. ;
		weights:long_name = "Ensemble weights" ;
		weights:comment = "No comments" ;
		weights:_FillValue = -9900. ;
		weights:valid_min = 0. ;
		weights:valid_max = 1. ;

// global attributes:
		:comment = "No comments" ;
		:Conventions = "CF-1.5 UW-1.0" ;
		:history = "No history" ;
		:institution = "NILU - Norwegian Institute for Air Research (http://www.nilu.no)" ;
		:references = "No references" ;
		:source = "No source" ;
		:title = "No title" ;
		:primary_variables = "no2_conc_grid_ctl no2_conc_grid_ens" ;
data:

 x = -14500, -13500, -12500, -11500, -10500, -9500, -8500, -7500, -6500,
    -5500, -4500, -3500, -2500, -1500, -500, 500, 1500, 2500, 3500, 4500,
    5500, 6500, 7500, 8500, 9500, 10500, 11500, 12500, 13500, 14500 ;

 y = -14500, -13500, -12500, -11500, -10500, -9500, -8500, -7500, -6500,
    -5500, -4500, -3500, -2500, -1500, -500, 500, 1500, 2500, 3500, 4500,
    5500, 6500, 7500, 8500, 9500, 10500, 11500, 12500, 13500, 14500 ;

 z = 1 ;

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19,
    20, 21, 22, 23, 24 ;

 no2_conc_grid_ctl =
  5.883742, 4.964289, 5.343208, 5.426654, 5.497732, 5.617154, 5.822791,
    6.085476, 6.551413, 7.475598, 9.228534, 11.34511, 12.99426, 16.53525,
    20.64528, 25.36003, 30.73264, 35.79173, 40.98288, 46.52135, 52.19265,
    56.94482, 60.4026, 62.61406, 63.61765, 61.39655, 59.59712, 62.09688,
    56.54461, 54.32262,
  4.59071, 3.909204, 4.201281, 4.69194, 4.936469, 5.117355, 5.450998,
    5.664864, 5.943838, 6.563833, 7.944495, 10.37015, 13.58713, 16.5691,
    20.35414, 25.83289, 30.86249, 35.99063, 41.70974, 47.88648, 53.35267,
    58.16707, 61.67268, 63.82231, 64.69511, 64.09298, 59.60417, 60.92033,
    56.78565, 54.94981,
  7.248794, 6.998601, 7.921134, 8.486769, 9.267927, 10.14715, 10.88618,
    11.54232, 11.99302, 12.36188, 12.88282, 14.00212, 15.96288, 18.83227,
    22.26036, 25.69117, 31.32148, 36.9812, 43.01134, 49.42927, 55.49656,
    60.42731, 63.82695, 65.409, 65.57798, 65.02164, 64.53706, 62.03141,
    55.92933, 54.88562,
  9.922905, 10.14669, 11.4794, 12.39308, 12.6625, 12.81061, 12.93595,
    13.04779, 13.36007, 14.02504, 15.14761, 16.60394, 18.60395, 21.40234,
    24.79404, 28.43181, 32.63522, 37.21527, 43.07146, 49.49315, 55.73454,
    60.69253, 63.64534, 65.63593, 65.91368, 65.8395, 65.76759, 64.78529,
    63.58326, 55.57288,
  12.5342, 12.60156, 13.03413, 12.99498, 13.06406, 13.06061, 13.11686,
    13.17702, 13.52216, 14.38081, 15.79214, 17.79613, 20.10247, 22.86383,
    26.06639, 29.80175, 34.04123, 38.76861, 44.25089, 50.69655, 56.32738,
    60.30507, 63.48089, 65.24516, 65.72262, 65.6589, 65.45322, 66.21934,
    65.81213, 63.8868,
  12.12335, 12.71982, 13.25724, 13.43924, 13.54796, 13.54546, 13.74328,
    13.87848, 13.9372, 14.42782, 15.69421, 17.76015, 20.57956, 23.47517,
    26.81104, 30.81075, 35.70746, 40.71364, 46.08905, 52.05994, 57.17648,
    60.86267, 63.88076, 65.16444, 65.42238, 65.1842, 64.70047, 65.22636,
    65.17465, 59.41511,
  12.37502, 12.67535, 13.24035, 13.43182, 13.69108, 13.94515, 14.33233,
    14.74863, 15.08075, 15.50035, 16.37879, 17.58301, 18.21667, 22.13759,
    25.68463, 29.87294, 34.65276, 40.22553, 45.78075, 52.13626, 57.47038,
    61.54484, 64.196, 65.53738, 65.59959, 64.95665, 64.79755, 64.89506,
    64.20908, 52.88522,
  14.1848, 13.08425, 13.56361, 13.62846, 13.78238, 14.21888, 14.57079,
    13.67422, 11.69121, 14.41622, 15.60628, 17.35281, 19.65482, 22.64098,
    26.193, 29.95635, 34.81673, 40.48651, 46.33178, 52.40357, 57.85375,
    61.94355, 64.55042, 65.67285, 65.5079, 65.26743, 65.39887, 64.90961,
    63.55021, 53.18229,
  16.9232, 15.07002, 14.91976, 14.61829, 14.42554, 14.34236, 13.46328,
    13.42105, 13.74318, 14.29393, 16.0461, 17.98164, 20.31268, 23.34734,
    26.8885, 30.11884, 34.79385, 40.9637, 47.342, 53.32038, 58.55437,
    62.61028, 64.88095, 65.49088, 65.20593, 65.56253, 65.47585, 64.43912,
    53.37814, 53.76642,
  21.7746, 19.58822, 18.27187, 17.17089, 16.66054, 15.71116, 13.95671,
    14.2232, 14.26684, 14.90268, 16.36649, 18.9205, 21.54687, 23.84576,
    26.62593, 30.58757, 35.34128, 40.81249, 46.96486, 53.44427, 59.26716,
    63.04467, 64.45132, 64.37296, 64.74198, 65.13624, 64.76041, 59.88474,
    53.06495, 52.83985,
  26.63352, 23.8249, 23.78424, 21.46133, 20.33435, 18.54521, 16.97405,
    16.00294, 15.83401, 16.62502, 17.54267, 19.41808, 21.37405, 24.19057,
    27.51903, 31.04685, 35.54198, 40.69891, 46.43068, 52.45237, 58.88805,
    62.84497, 64.14728, 64.33866, 64.74864, 64.46625, 61.46327, 53.45512,
    54.00876, 52.93948,
  27.30437, 24.70839, 27.33698, 27.52127, 26.32023, 22.79061, 19.65536,
    16.74692, 15.6199, 16.33771, 17.62616, 19.55305, 22.56422, 25.09051,
    27.96906, 32.12367, 35.9793, 40.98378, 46.70205, 52.40247, 58.03683,
    62.4975, 63.86574, 64.68283, 64.93655, 64.10212, 53.72129, 57.71857,
    54.54689, 53.59676,
  17.69748, 18.81306, 21.01472, 23.86465, 25.94342, 25.55343, 19.5307,
    14.43942, 17.98577, 17.01037, 18.62759, 19.98468, 22.35567, 24.98332,
    28.15253, 31.38074, 36.12353, 41.32821, 47.07075, 52.92445, 58.22942,
    61.91414, 63.6117, 63.37764, 63.21084, 62.02723, 54.45757, 55.96704,
    55.4805, 54.3599,
  13.96198, 12.64386, 12.82304, 13.05641, 13.62405, 14.39063, 15.31632,
    16.51217, 15.56489, 16.8012, 18.76303, 21.04775, 23.13984, 25.34055,
    28.59778, 31.90468, 35.63426, 41.75359, 47.91163, 53.57299, 58.00996,
    61.30392, 61.42176, 57.0647, 54.13472, 54.41312, 53.89153, 53.47883,
    53.69308, 53.73604,
  14.80429, 11.35051, 14.17216, 14.15507, 14.40264, 14.54152, 14.84269,
    15.02591, 15.5501, 17.00052, 18.88947, 21.1168, 23.47238, 26.16829,
    28.56116, 31.63985, 36.31792, 40.36988, 46.90042, 53.18296, 55.71748,
    59.02044, 57.07051, 55.24336, 55.60468, 54.81219, 54.1027, 53.61647,
    53.17145, 53.06683,
  9.873219, 10.90184, 12.65371, 13.79382, 14.20805, 14.73239, 15.35361,
    15.70504, 16.36293, 18.16138, 20.68384, 22.84251, 25.10741, 26.87732,
    29.38061, 32.63404, 36.01141, 40.34125, 44.92809, 49.90028, 51.39642,
    55.31063, 55.46692, 55.39748, 55.36237, 54.77618, 54.02326, 53.61515,
    53.24664, 53.10964,
  7.219785, 5.595117, 7.13706, 8.640588, 10.43177, 12.76819, 14.17335,
    14.9413, 16.19319, 18.20708, 20.58299, 23.58203, 27.07339, 29.36787,
    31.81454, 34.51089, 37.65513, 42.12624, 47.68143, 51.3913, 51.82205,
    55.43442, 55.79317, 55.44896, 55.30649, 54.92293, 53.97525, 53.19198,
    52.97479, 52.98631,
  10.39959, 7.227608, 6.212149, 6.50093, 7.710369, 8.86208, 10.24349,
    11.81669, 14.18129, 16.06364, 18.71134, 22.13064, 25.44047, 29.99675,
    33.7595, 36.74979, 40.07243, 45.07722, 51.11308, 56.1602, 54.92405,
    55.88823, 56.00541, 55.92464, 55.22741, 54.75513, 54.08841, 53.07667,
    52.82054, 52.86615,
  23.8078, 16.14485, 9.081383, 4.16374, 6.090626, 6.253955, 7.258926,
    8.351885, 9.510268, 11.65442, 15.14532, 18.04436, 20.30593, 26.49682,
    32.10813, 36.56562, 41.57413, 47.91143, 54.78819, 60.01239, 62.55959,
    59.81793, 57.5056, 57.34682, 55.99229, 55.21619, 54.44096, 53.27673,
    52.78887, 52.88083,
  23.42601, 16.41229, 9.401606, 4.596685, 6.022668, 6.261339, 7.17676,
    8.310963, 10.16568, 13.06719, 15.43149, 15.63903, 18.73225, 21.54271,
    25.41957, 30.41687, 37.24792, 45.6711, 52.73322, 58.48302, 62.4933,
    62.59989, 59.61031, 58.64321, 57.17355, 55.6868, 54.67691, 53.4545,
    52.7585, 52.90039,
  24.51663, 18.59818, 11.36408, 6.748722, 7.66969, 7.578695, 8.261253,
    9.202785, 10.90752, 13.01413, 14.06653, 15.16191, 19.38181, 22.40535,
    25.62338, 29.96549, 35.52126, 42.28676, 49.2677, 55.06973, 59.52965,
    62.36836, 61.92377, 60.19802, 58.28825, 56.19801, 54.69009, 53.45536,
    52.78088, 52.90583,
  25.20035, 21.35663, 15.01315, 11.26674, 12.7185, 12.17463, 12.66978,
    13.06605, 14.62867, 15.96196, 16.0278, 17.52586, 21.00344, 24.2227,
    27.50082, 31.83625, 36.94009, 42.8319, 48.82259, 53.81068, 57.82055,
    60.30282, 61.88569, 61.83137, 60.05999, 57.11857, 55.16679, 53.92423,
    52.8901, 52.88246,
  25.64075, 22.32646, 18.01783, 15.02031, 17.70362, 18.5392, 19.19979,
    19.22233, 20.08348, 20.73996, 21.33334, 24.38845, 27.63299, 30.76249,
    33.62913, 37.58646, 42.19489, 46.71119, 51.46165, 55.43668, 58.56087,
    60.48229, 61.1334, 61.42413, 61.73009, 59.21924, 56.34901, 54.84444,
    53.66804, 53.01262,
  25.61953, 22.23292, 18.95841, 17.29291, 18.54148, 19.10852, 20.35045,
    21.88209, 23.70866, 25.0326, 27.03034, 30.60055, 34.61942, 38.14453,
    41.15078, 44.87738, 49.14297, 53.58028, 57.06005, 60.47861, 62.75799,
    63.41985, 62.74937, 62.17194, 62.51088, 62.14661, 59.64099, 56.21656,
    54.83282, 53.77882,
  25.40796, 21.2502, 17.80196, 14.81898, 16.78609, 17.52773, 18.84142,
    20.79207, 22.83847, 24.27811, 26.28782, 29.95529, 34.29748, 38.11113,
    41.12055, 45.00898, 49.28408, 53.97094, 58.83229, 62.79018, 65.21492,
    65.68035, 63.90536, 62.31511, 62.41687, 62.22562, 61.32932, 57.98138,
    55.5217, 54.52943,
  27.25072, 23.27057, 19.78855, 17.39992, 17.97907, 18.57905, 20.27608,
    22.34326, 24.05668, 25.45224, 27.9048, 31.33662, 35.48065, 38.92867,
    41.66696, 45.27874, 49.28631, 53.69078, 58.52177, 63.26844, 66.48228,
    67.53506, 66.01924, 64.24088, 63.8571, 62.83379, 62.01669, 59.07139,
    55.08469, 54.03268,
  35.6475, 32.10685, 28.71725, 26.47991, 26.88938, 26.3118, 28.36579,
    29.8306, 30.26041, 31.42297, 34.55059, 38.33418, 41.91167, 44.79679,
    46.9156, 49.6423, 52.23276, 55.48059, 59.42588, 63.37962, 66.16835,
    67.75281, 67.37491, 66.17617, 65.7543, 64.9575, 64.6252, 62.39565,
    56.8582, 53.65231,
  48.6854, 47.0442, 44.2873, 42.8579, 43.79852, 44.16705, 44.19046, 43.51111,
    42.50537, 43.387, 44.69755, 47.11941, 50.3853, 52.87177, 53.90959,
    55.14336, 55.94797, 57.39343, 59.99869, 63.06133, 64.27831, 64.19556,
    63.16653, 62.36388, 62.64981, 62.45007, 62.10195, 61.95482, 59.93761,
    55.14679,
  53.94149, 54.59158, 55.85206, 56.51167, 57.37472, 58.35294, 58.55539,
    54.45732, 53.1251, 53.58015, 53.30247, 53.52778, 54.19484, 55.02066,
    55.52387, 55.87267, 55.80025, 55.99661, 56.42194, 56.9221, 57.86377,
    58.90435, 59.02439, 58.41271, 58.62147, 58.60619, 58.04326, 56.58253,
    56.01933, 55.15231,
  57.13857, 57.73228, 58.06318, 58.05644, 59.28595, 61.71721, 62.00758,
    58.48709, 56.28851, 57.10241, 57.56494, 58.1425, 58.19043, 57.79145,
    57.27106, 56.82783, 55.71459, 54.46612, 54.3838, 54.49223, 54.29781,
    55.03545, 55.88245, 56.26332, 56.18774, 56.44104, 56.13518, 54.95704,
    53.85836, 53.08151,
  26.32195, 28.39637, 30.86953, 33.49986, 36.34968, 39.41561, 42.5379,
    45.68922, 48.94297, 52.23912, 55.55793, 58.55124, 60.74559, 62.47725,
    63.64361, 64.31554, 64.64057, 64.82305, 64.93568, 65.02431, 64.89962,
    64.47733, 64.06298, 63.74698, 63.27929, 62.48074, 55.46485, 58.1342,
    54.18584, 51.62521,
  25.54156, 27.57197, 30.29865, 33.12555, 36.19661, 39.48579, 43.00047,
    46.40277, 49.77276, 53.15023, 56.44667, 59.59335, 62.05659, 63.64996,
    64.46265, 64.85717, 64.97762, 65.06114, 65.1627, 65.438, 65.66352,
    65.69538, 65.58854, 65.41722, 65.12701, 63.87126, 62.19883, 56.89033,
    53.56446, 51.94366,
  26.49522, 28.40215, 31.06346, 33.77855, 36.66869, 39.74959, 43.26157,
    46.99924, 50.61823, 54.05937, 57.14748, 60.06356, 62.54142, 64.27589,
    65.18645, 65.31932, 65.2205, 65.17213, 65.17397, 65.20673, 65.5928,
    66.0714, 66.11716, 65.91725, 65.41304, 64.951, 64.28798, 62.5515,
    54.19318, 51.62819,
  26.89033, 29.07411, 31.96473, 34.63583, 37.38411, 40.17265, 43.32393,
    46.99594, 50.72496, 54.50309, 57.81824, 60.67699, 63.15678, 64.81903,
    65.78314, 66.10425, 65.80836, 65.5362, 65.60097, 65.5663, 65.70992,
    65.57636, 64.82198, 65.02841, 64.66375, 64.91461, 65.22162, 64.4421,
    62.66006, 54.52505,
  27.39697, 29.72588, 32.78268, 35.96497, 38.59081, 41.15557, 43.81313,
    47.2177, 50.5288, 54.2332, 57.69999, 60.87417, 63.76014, 65.57325,
    66.50533, 66.89861, 66.67197, 66.20085, 66.04906, 65.98981, 65.54056,
    64.67014, 64.56243, 64.57603, 64.39697, 64.24498, 64.30313, 65.38677,
    64.98656, 62.55223,
  28.26976, 30.16733, 33.22097, 36.40108, 39.57649, 42.21046, 44.66718,
    48.19107, 51.18317, 54.1033, 57.27514, 60.55339, 63.728, 65.62126,
    66.85735, 67.51149, 67.24005, 66.7958, 66.18807, 65.92648, 65.3391,
    64.42715, 64.7761, 64.76933, 64.5081, 64.11785, 63.72606, 64.295,
    64.25084, 56.8594,
  31.40828, 32.06876, 34.23016, 36.84999, 39.85476, 42.77045, 45.50473,
    48.85038, 52.19762, 55.05081, 57.82937, 60.07606, 61.54239, 63.61354,
    64.95271, 65.79875, 66.20486, 65.82112, 65.00177, 64.85339, 64.62834,
    64.52828, 64.69029, 64.9002, 64.62935, 64.17639, 64.06433, 64.00343,
    63.18209, 50.16885,
  36.68778, 36.38324, 37.26472, 38.71168, 40.91144, 43.91642, 46.82381,
    48.2878, 50.68326, 53.69422, 56.40186, 58.96917, 61.27497, 63.31631,
    64.79969, 65.54571, 66.16996, 66.38718, 65.87499, 65.1723, 64.72418,
    64.5475, 64.57025, 64.60274, 64.29213, 64.29124, 64.42776, 63.75282,
    62.07674, 50.4953,
  42.50343, 42.86539, 42.72434, 42.94631, 43.80785, 45.60265, 46.68948,
    49.08482, 52.01757, 54.69712, 57.15117, 59.36504, 61.19577, 63.07761,
    64.67322, 65.14552, 65.77427, 66.60606, 66.91232, 66.30061, 65.55784,
    64.91251, 64.4489, 63.95583, 63.7194, 64.26557, 64.23694, 63.02283,
    50.32836, 51.03104,
  45.54002, 48.34453, 49.23274, 49.03627, 48.68483, 48.54872, 48.36039,
    50.49408, 52.98457, 55.80845, 57.98517, 60.02913, 61.50135, 62.60313,
    63.41371, 64.43441, 65.04243, 65.55288, 65.98151, 66.06835, 66.14948,
    65.21802, 64.18037, 63.26911, 63.40537, 63.66018, 63.23866, 57.42121,
    50.56318, 50.26687,
  44.1024, 47.17902, 51.65185, 53.79406, 54.1587, 53.00584, 52.44597,
    52.95064, 54.29271, 57.20134, 59.01999, 60.25147, 61.45216, 62.4181,
    63.14435, 63.78362, 64.26437, 64.50961, 64.78033, 64.91776, 65.58309,
    65.07374, 63.76572, 63.42927, 63.84787, 63.3275, 60.66906, 51.79583,
    51.6624, 50.55094,
  40.38974, 40.62097, 47.89691, 53.63884, 58.45015, 57.59234, 55.27719,
    53.62546, 55.48582, 57.27234, 59.53749, 61.02785, 62.7731, 63.61884,
    63.84853, 63.99577, 64.48349, 64.72112, 64.71497, 64.54523, 64.9998,
    64.81435, 63.46838, 63.20876, 63.54166, 62.88597, 50.69913, 56.26461,
    52.58034, 51.3895,
  34.45702, 37.16591, 40.12017, 46.01087, 52.40127, 57.21019, 55.49479,
    52.49266, 58.25724, 59.01358, 61.348, 62.70934, 64.23479, 65.3399,
    65.49723, 64.23989, 64.69238, 65.19176, 65.23018, 64.71075, 64.72763,
    64.41058, 63.53138, 60.85248, 58.93715, 60.29039, 51.26732, 52.57795,
    53.0231, 52.11128,
  32.48871, 34.73455, 36.61579, 39.3309, 42.32029, 45.69027, 50.41014,
    55.27252, 56.64538, 59.56109, 62.27788, 64.45454, 65.60512, 66.48157,
    66.63222, 65.70441, 64.90005, 65.20869, 65.64873, 64.86847, 63.91064,
    63.31743, 61.4445, 55.65688, 51.17601, 51.3297, 51.38934, 50.53649,
    50.72923, 51.08976,
  30.62918, 29.78183, 35.75975, 38.99873, 42.34248, 45.74797, 48.67188,
    52.10448, 56.24026, 59.55516, 61.94947, 63.88294, 65.66982, 67.01015,
    67.30505, 67.34953, 66.33867, 65.08515, 64.56281, 64.20516, 60.58063,
    60.38355, 56.18478, 52.89112, 53.30016, 52.11507, 51.49426, 51.02335,
    50.47031, 50.39288,
  26.16108, 28.71323, 31.68517, 35.82912, 40.09167, 43.70455, 46.98085,
    50.42199, 54.17956, 58.15782, 61.32863, 63.64425, 65.66732, 67.39745,
    68.05708, 68.07531, 67.81328, 66.51816, 64.97314, 61.29711, 57.66827,
    57.2005, 54.81155, 53.26023, 52.78441, 52.04896, 51.18523, 50.81309,
    50.55823, 50.49673,
  30.06777, 28.76213, 31.93294, 34.91405, 38.40325, 42.10611, 46.47615,
    49.46418, 52.69479, 56.2701, 59.5248, 62.73822, 65.58553, 67.10249,
    68.09168, 68.92403, 69.37775, 68.97482, 67.68057, 65.84844, 59.44137,
    57.86348, 55.66923, 53.86373, 53.11073, 52.3774, 51.23965, 50.49348,
    50.34087, 50.36295,
  40.26164, 36.29704, 34.90982, 36.35675, 40.25679, 43.42276, 47.13813,
    50.68885, 53.55054, 56.39506, 59.3933, 62.36061, 64.36369, 65.85339,
    66.73769, 67.9621, 69.38531, 70.36554, 70.399, 68.96164, 65.88673,
    59.5316, 56.55768, 55.17062, 53.29605, 52.6293, 51.63862, 50.51403,
    50.28896, 50.28436,
  50.27216, 46.6272, 42.31796, 37.16735, 42.0353, 44.73307, 48.42007,
    51.88935, 55.47208, 58.69918, 61.27591, 63.30339, 63.23682, 63.38673,
    63.67083, 65.5792, 67.67566, 69.29895, 70.25424, 70.35391, 68.86745,
    64.67379, 58.39419, 57.22223, 54.7353, 53.53791, 52.45162, 50.81499,
    50.25414, 50.31215,
  49.98399, 47.20474, 43.76025, 40.78366, 44.8838, 47.332, 51.04577,
    54.74586, 58.16003, 61.17732, 63.4836, 65.09465, 66.66003, 66.97263,
    65.28389, 64.24108, 64.69789, 66.61615, 67.76351, 67.73814, 67.61839,
    66.55026, 61.15645, 58.5395, 56.34575, 54.34702, 52.93164, 51.09134,
    50.13005, 50.32421,
  51.41594, 48.68894, 45.34512, 44.20398, 47.96408, 50.54058, 53.79267,
    57.13945, 60.65248, 63.61625, 65.90346, 67.38584, 68.89587, 69.63257,
    69.58329, 68.77944, 67.89446, 67.63426, 67.1697, 65.69092, 64.98389,
    64.9267, 63.21612, 60.26765, 57.83756, 55.22976, 53.1363, 51.27039,
    50.17722, 50.29074,
  54.74319, 52.05514, 48.52501, 47.35733, 51.15362, 53.67402, 56.96374,
    60.04397, 63.42273, 66.73827, 69.29752, 71.19158, 72.49226, 72.92081,
    72.7149, 72.15528, 71.2761, 70.15755, 69.03141, 67.04601, 65.33289,
    63.63001, 63.21078, 61.64175, 59.73863, 56.35162, 53.87782, 52.10767,
    50.60505, 50.32993,
  61.25042, 58.47228, 54.53007, 52.89367, 56.13809, 58.46863, 61.49236,
    64.34846, 67.24219, 70.06226, 72.90993, 75.77758, 77.71684, 78.0572,
    77.41789, 76.67329, 75.5462, 74.10522, 72.60812, 70.80087, 68.30486,
    65.97838, 63.68814, 62.21605, 61.76838, 58.88145, 55.22875, 53.25972,
    51.76306, 50.64307,
  69.20071, 65.92104, 61.78536, 59.8088, 61.94831, 63.3198, 65.73111,
    68.54162, 71.54849, 73.51946, 75.70938, 79.13476, 82.28674, 83.41745,
    82.43775, 81.66219, 80.37843, 78.65395, 76.74957, 75.21064, 73.71432,
    70.36469, 66.36801, 63.69684, 63.11646, 61.70776, 58.62987, 54.60664,
    52.97832, 51.60237,
  75.48962, 71.65627, 66.61379, 63.74545, 65.01375, 65.54831, 67.10264,
    69.53745, 72.28286, 73.5099, 74.99456, 77.60227, 80.5438, 81.91639,
    81.03331, 80.63384, 79.65504, 78.46567, 77.16338, 75.87045, 74.57363,
    72.17223, 67.33808, 64.22171, 63.58058, 62.34664, 60.40053, 56.26242,
    53.16819, 52.18768,
  78.34026, 73.95398, 68.88648, 65.55232, 65.52935, 64.99583, 67.27913,
    69.16975, 70.78522, 71.19975, 72.52689, 74.85516, 77.92771, 78.96007,
    78.16717, 77.98851, 77.36433, 76.41665, 75.38326, 74.64208, 73.33362,
    71.10536, 67.2725, 64.42483, 63.97662, 62.84865, 61.57186, 57.9339,
    53.15634, 51.60944,
  76.67091, 73.1258, 68.38963, 65.06921, 65.09248, 63.32303, 64.11791,
    65.39435, 65.67062, 65.04703, 66.31236, 69.15531, 73.31841, 74.92999,
    74.20624, 73.73901, 72.88653, 72.08736, 71.24966, 70.78586, 69.96158,
    68.44622, 65.54892, 63.32589, 63.06023, 62.5658, 62.04759, 60.03755,
    55.09871, 51.58838,
  70.81985, 69.09328, 65.90504, 63.90758, 64.73823, 63.96408, 62.67867,
    61.8185, 60.85789, 60.59913, 60.24672, 61.56745, 64.71053, 66.71094,
    66.25034, 65.76791, 64.86174, 64.0207, 63.856, 64.63331, 64.56799,
    63.436, 60.99949, 59.44199, 59.62309, 59.18034, 58.29462, 57.66132,
    56.49603, 52.71521,
  56.74456, 57.59261, 58.99742, 60.27051, 61.42245, 63.17837, 61.23394,
    57.53094, 56.34059, 56.81397, 56.2406, 55.80711, 55.91445, 56.53045,
    56.65422, 56.40686, 55.80711, 55.20919, 54.70458, 54.56804, 55.12868,
    56.20812, 56.56524, 55.91032, 56.19289, 56.14516, 55.32659, 53.43466,
    52.53767, 52.19289,
  54.09917, 54.43099, 54.8211, 54.8234, 55.48502, 57.03102, 57.7861,
    55.12793, 53.40697, 54.1084, 54.43875, 54.55325, 54.3008, 54.03064,
    53.8833, 53.6216, 52.74176, 51.65251, 51.44669, 51.44159, 51.16365,
    51.72047, 52.69196, 53.22492, 53.20388, 53.42119, 53.20483, 52.11079,
    51.05979, 50.45716,
  58.99273, 60.61912, 61.56118, 62.54097, 63.18652, 63.63482, 63.84388,
    63.96794, 63.96114, 63.8157, 63.64489, 63.53851, 63.34473, 63.24617,
    63.11407, 62.99908, 63.02084, 63.26271, 63.46997, 63.53006, 63.28553,
    62.88264, 62.56121, 62.19721, 61.83627, 54.7692, 49.73812, 51.95679,
    49.28982, 47.44821,
  58.83477, 60.45273, 61.4419, 62.49816, 63.15544, 63.65, 63.99109, 64.16876,
    64.2427, 64.29456, 64.12485, 64.00149, 63.92965, 63.66299, 63.34454,
    63.14714, 63.06728, 63.25747, 63.51522, 63.76989, 63.88236, 64.0028,
    63.88961, 63.78935, 63.33163, 61.93058, 53.09292, 50.01264, 48.74421,
    47.60617,
  58.91188, 60.46044, 61.44778, 62.44239, 63.12868, 63.6707, 63.9487,
    64.1256, 64.22794, 64.26988, 64.30832, 64.23344, 64.11082, 64.02854,
    63.80688, 63.49546, 63.32999, 63.27212, 63.29753, 63.46498, 63.89349,
    64.26723, 64.51376, 64.47127, 63.88442, 63.11087, 62.12548, 56.37332,
    48.73529, 47.53164,
  59.0666, 60.53911, 61.46357, 62.44384, 63.20778, 63.86753, 64.20644,
    64.24414, 64.30795, 64.28577, 64.33296, 64.59634, 64.69083, 64.42049,
    64.26755, 64.18506, 63.89071, 63.57169, 63.52768, 63.56797, 63.81996,
    63.77797, 63.20567, 63.57248, 63.37999, 63.43342, 63.28931, 62.5386,
    60.90261, 49.81509,
  59.32707, 60.6915, 61.53933, 62.35302, 63.02967, 63.74174, 64.37505,
    64.52739, 64.37766, 64.25493, 64.31773, 64.92861, 65.47633, 65.18948,
    64.9859, 64.79769, 64.58039, 64.19145, 64.03495, 63.89548, 63.42261,
    62.84532, 62.33656, 63.10826, 63.12273, 62.97507, 63.00948, 63.81895,
    63.59995, 60.14583,
  59.94938, 61.06391, 61.9815, 62.71337, 63.10825, 63.65379, 64.47419,
    65.00019, 64.94043, 64.73864, 64.82631, 65.2428, 65.90161, 65.68551,
    65.51241, 65.36503, 64.77846, 64.57341, 64.4265, 64.04948, 63.40824,
    60.96272, 63.0204, 63.12844, 63.01127, 62.83476, 62.5793, 62.91398,
    62.90403, 52.53861,
  61.84982, 62.01446, 62.76665, 63.27027, 63.61055, 64.084, 64.71255,
    64.89105, 64.94902, 64.93957, 65.00095, 64.65079, 63.87796, 64.14643,
    64.16896, 64.12714, 64.08943, 63.59766, 63.03294, 62.99841, 62.71292,
    62.62312, 62.84687, 63.16108, 63.09216, 62.87912, 62.8882, 62.8844,
    62.12691, 46.45356,
  65.90823, 64.64047, 64.43394, 64.44605, 64.50874, 65.00803, 65.30882,
    63.89402, 62.95273, 62.97055, 63.12128, 63.23998, 63.50694, 63.91435,
    64.22456, 64.31598, 64.34823, 64.21466, 63.69798, 63.18126, 62.82588,
    62.67875, 62.75117, 62.8842, 62.82616, 63.00003, 63.15757, 62.54477,
    59.29828, 46.72211,
  71.43134, 70.25322, 68.2494, 67.04137, 66.28838, 65.8057, 64.44878,
    64.32702, 63.88993, 63.39457, 63.20545, 63.16564, 63.03621, 63.39071,
    63.85721, 63.87615, 64.3046, 64.7917, 64.83825, 64.15795, 63.61903,
    63.16401, 62.82813, 62.43147, 62.26576, 62.80814, 62.97716, 62.00307,
    46.63613, 47.14249,
  74.54456, 76.01109, 74.47547, 72.26646, 70.12727, 67.85751, 65.37211,
    65.24444, 64.85873, 64.45671, 63.71859, 63.2162, 62.79732, 62.63943,
    62.36097, 62.26917, 62.63955, 63.83066, 64.2791, 64.20501, 64.13409,
    63.49207, 62.78352, 62.09308, 62.17436, 62.21528, 61.98483, 53.04245,
    46.69509, 46.69498,
  72.61015, 75.31149, 78.46147, 77.98033, 76.01496, 71.72469, 68.55814,
    66.64463, 65.62534, 65.84274, 64.53073, 63.13266, 62.6273, 62.34212,
    62.15729, 62.10856, 60.72142, 59.58612, 59.76798, 61.24554, 63.67282,
    63.30425, 62.39029, 62.34227, 62.96021, 62.59674, 56.15246, 47.51489,
    47.73571, 46.81566,
  68.57148, 68.75275, 74.1528, 78.1844, 79.39154, 75.95925, 71.3905,
    67.74648, 66.50908, 66.05348, 65.29458, 64.33368, 64.00869, 63.61049,
    62.8858, 62.49839, 62.69586, 62.84123, 61.12144, 60.04893, 62.17859,
    62.82301, 61.42433, 61.94366, 62.48124, 62.18869, 47.19526, 52.2248,
    48.44685, 47.48691,
  62.69732, 64.49674, 66.09728, 69.5303, 72.96391, 74.54807, 70.13905,
    66.52438, 68.77477, 67.48044, 66.86735, 65.90947, 65.7207, 65.4132,
    64.51657, 62.71196, 62.94947, 63.28822, 63.28295, 62.90216, 63.12469,
    62.97707, 61.78868, 55.67397, 54.40425, 56.10628, 47.57326, 49.14901,
    49.12132, 48.14334,
  62.94706, 63.79455, 63.73693, 62.92904, 62.24274, 64.4846, 66.61392,
    68.05413, 66.51142, 67.39615, 67.6768, 67.01656, 66.5779, 66.28987,
    65.27167, 63.79776, 63.07839, 63.38419, 63.81198, 63.23412, 62.60152,
    62.08929, 55.06553, 50.26347, 47.01863, 47.29499, 47.53803, 46.86694,
    47.12562, 47.34743,
  63.30683, 63.36695, 64.95009, 65.03533, 65.00662, 65.25911, 65.79366,
    65.97727, 65.89526, 65.7983, 65.99385, 65.96815, 66.24542, 66.15253,
    65.47289, 65.0574, 63.86603, 63.24125, 63.1247, 62.05961, 55.54506,
    55.14156, 51.54345, 48.26695, 48.79066, 48.09802, 47.6225, 47.22524,
    46.78013, 46.74929,
  61.27607, 63.54976, 64.41871, 65.08394, 65.31263, 65.66931, 66.11597,
    66.16689, 65.67509, 65.22459, 65.38597, 65.77763, 66.32122, 66.96931,
    66.418, 65.58017, 65.19653, 64.25597, 59.05282, 56.24641, 53.33377,
    52.21341, 49.97488, 48.64044, 48.42502, 47.99948, 47.42266, 47.06848,
    46.83742, 46.84087,
  64.98389, 64.56703, 65.2938, 65.73668, 65.53836, 65.5983, 66.03209,
    66.66262, 66.24703, 65.53658, 65.134, 65.68341, 66.72715, 67.02293,
    66.93155, 67.06305, 67.08855, 66.67413, 65.24268, 60.42118, 54.58601,
    52.9625, 50.84876, 49.24316, 48.89399, 48.35628, 47.42813, 46.81373,
    46.70806, 46.72623,
  71.96576, 70.12035, 67.32001, 66.91241, 67.61699, 67.36596, 67.45039,
    67.41502, 67.41074, 66.31326, 66.21727, 66.19176, 66.05421, 65.84758,
    65.79841, 66.64999, 67.81297, 68.46161, 68.19569, 66.65241, 60.08804,
    54.59923, 51.92299, 50.63725, 49.26643, 48.72559, 47.73595, 46.84416,
    46.62959, 46.65303,
  81.3079, 77.27425, 72.35072, 66.95946, 69.24029, 68.60318, 68.69923,
    68.59464, 67.68616, 67.61959, 67.64951, 66.8713, 64.06648, 61.99721,
    60.68012, 61.9879, 65.87712, 67.68375, 68.37181, 68.35953, 66.86632,
    59.3763, 53.90604, 52.75148, 50.63043, 49.61026, 48.56308, 47.06979,
    46.56023, 46.65335,
  80.66859, 77.28825, 72.55075, 68.35941, 70.44502, 70.49426, 70.46449,
    70.18102, 70.16288, 69.85267, 69.43987, 68.95763, 68.5452, 65.58026,
    62.49611, 60.8905, 60.99, 62.48818, 63.24579, 63.70645, 63.44025,
    60.64824, 56.20382, 54.05409, 52.00499, 50.31384, 49.02724, 47.34479,
    46.47858, 46.67783,
  80.39993, 77.24596, 72.36029, 68.75802, 70.92812, 71.01414, 71.84628,
    72.27644, 72.52014, 72.12904, 70.7272, 69.26598, 69.51772, 68.78642,
    66.87959, 65.60505, 64.74699, 64.25154, 63.38989, 61.35248, 59.68482,
    58.90779, 57.57861, 55.22824, 53.39695, 51.17213, 49.25268, 47.46215,
    46.49853, 46.64333,
  78.81881, 76.3017, 71.46362, 68.11389, 70.88901, 71.42703, 72.49573,
    73.22865, 74.06618, 74.54298, 74.25061, 73.16388, 72.41711, 71.30345,
    70.21146, 69.06589, 67.61997, 66.58965, 65.38847, 63.11814, 60.39046,
    57.98157, 57.95401, 56.07484, 54.6195, 52.20302, 50.08601, 48.15864,
    46.75648, 46.64638,
  77.92939, 75.21868, 70.22502, 66.87189, 69.75492, 70.84918, 72.10115,
    73.07625, 74.59246, 75.96823, 76.75008, 76.8734, 76.58264, 76.13665,
    75.28319, 74.39993, 73.24516, 71.2784, 69.19566, 66.47393, 63.33215,
    60.49627, 58.59526, 56.7981, 56.27824, 54.13087, 51.19721, 49.1706,
    47.64143, 46.87094,
  76.98052, 73.99052, 69.1778, 66.1955, 68.02755, 69.08877, 70.65472,
    72.55482, 74.69102, 76.13597, 77.26913, 79.006, 80.67355, 81.21273,
    80.14568, 79.37634, 77.91215, 76.23412, 74.39162, 71.56659, 68.88776,
    65.04192, 61.1142, 58.78173, 57.98057, 56.75744, 54.00548, 50.39775,
    48.76707, 47.61811,
  76.57349, 72.94313, 66.93142, 62.48405, 63.58941, 63.93969, 66.52797,
    69.7989, 72.80685, 73.72358, 74.51743, 76.28649, 78.9332, 80.0098,
    79.20049, 78.55952, 77.70691, 76.43222, 74.48882, 72.32039, 69.85645,
    66.63694, 62.3369, 59.36237, 58.74559, 57.24899, 55.33817, 51.74353,
    49.05864, 48.21722,
  76.01103, 72.29289, 66.53738, 61.46936, 61.34103, 60.7903, 62.7642,
    65.94393, 68.48134, 68.74431, 70.65054, 73.23837, 76.59114, 77.71593,
    76.55061, 76.10475, 74.67368, 73.44886, 71.98904, 70.81324, 68.985,
    66.3405, 62.59447, 59.8172, 59.26434, 57.73126, 56.13649, 53.04555,
    49.19369, 47.79087,
  73.77109, 70.95072, 64.89207, 60.26355, 60.44655, 58.99968, 59.59968,
    60.98069, 62.13649, 62.16152, 63.81998, 66.57539, 70.15773, 71.77969,
    70.98554, 70.09617, 69.11942, 67.74037, 67.56355, 67.27053, 66.38676,
    64.24622, 61.23448, 59.00227, 58.68431, 57.75036, 56.82928, 54.64824,
    50.69788, 47.79028,
  66.83418, 65.64572, 61.26554, 58.54013, 59.6647, 59.05951, 57.84234,
    57.30264, 56.93185, 56.74202, 56.92121, 58.32399, 61.15763, 63.01555,
    62.74211, 62.30353, 61.03873, 60.09299, 59.76657, 60.75104, 60.64718,
    59.61537, 57.22931, 55.57049, 55.72415, 55.03988, 54.11287, 53.20959,
    51.63136, 48.62328,
  52.29277, 53.32224, 54.48293, 55.30769, 56.33781, 57.74255, 56.16731,
    53.31594, 52.36998, 52.56065, 52.05969, 51.68238, 51.68433, 52.301,
    52.3829, 52.30188, 51.67092, 51.03308, 50.65427, 50.73912, 51.44331,
    52.39207, 52.79124, 52.17841, 52.1992, 52.18477, 51.41748, 49.81123,
    48.73994, 48.19281,
  49.65837, 50.06335, 50.56483, 50.58648, 51.21404, 52.60664, 52.99527,
    50.9696, 49.66304, 50.08705, 50.25576, 50.33722, 50.07931, 49.75881,
    49.61612, 49.42657, 48.71093, 47.8549, 47.66327, 47.65497, 47.53751,
    48.10098, 49.02553, 49.51527, 49.39439, 49.55245, 49.40165, 48.43999,
    47.47852, 46.86683,
  62.34592, 62.32872, 62.35643, 62.39123, 62.35184, 62.30035, 62.23705,
    61.82101, 60.94782, 60.24479, 59.89061, 59.82495, 59.70879, 60.54284,
    61.57648, 61.52942, 61.31005, 60.90985, 60.39878, 59.8817, 59.33674,
    58.75425, 56.30867, 54.51578, 52.21407, 48.50423, 45.81991, 47.36668,
    44.99749, 43.49381,
  62.64791, 62.73936, 62.70752, 62.72621, 62.69003, 62.63553, 62.58706,
    62.52792, 62.45068, 62.44021, 62.35231, 61.52407, 60.90967, 60.23229,
    60.19175, 61.30002, 61.3516, 61.17032, 60.96764, 60.75607, 60.46767,
    60.12526, 59.77248, 59.59562, 59.24296, 56.46268, 46.83749, 45.54879,
    44.69093, 43.64466,
  62.51096, 62.73236, 62.81153, 62.82334, 62.76603, 62.72168, 62.66064,
    62.58104, 62.53627, 62.50202, 62.46738, 62.45541, 62.30106, 62.14774,
    61.83683, 60.47123, 59.69016, 60.46129, 60.66764, 60.68728, 60.82327,
    60.92467, 60.86478, 60.61196, 59.91202, 58.8308, 58.11121, 48.86197,
    44.18914, 43.63903,
  62.44256, 62.66275, 62.83454, 62.96295, 63.01484, 63.07957, 63.00377,
    62.88665, 62.71206, 62.47709, 62.48372, 62.80302, 62.92252, 62.6467,
    62.40519, 62.02781, 61.3623, 60.69424, 60.42448, 60.46509, 60.62084,
    60.3554, 59.75237, 59.88795, 59.48848, 59.62163, 59.14415, 58.60843,
    53.26189, 45.16777,
  62.38734, 62.48444, 62.63798, 62.74805, 62.8188, 63.1339, 63.45832,
    63.34012, 63.0275, 62.60711, 62.49487, 63.08176, 63.63404, 63.35146,
    63.02103, 62.79724, 62.2692, 61.5284, 60.96095, 60.38846, 59.95313,
    57.8085, 54.9564, 57.059, 58.98971, 59.03974, 59.13326, 60.00146,
    60.02401, 54.69224,
  62.53683, 62.5606, 62.61914, 62.60093, 62.55066, 63.00255, 63.88382,
    64.25309, 64.05507, 63.59842, 63.3915, 63.75352, 64.28346, 63.81445,
    63.50825, 63.23818, 62.30818, 61.87815, 61.56681, 60.9658, 60.25692,
    54.86007, 58.31305, 57.60064, 57.50447, 57.04949, 57.53809, 59.04397,
    59.11611, 48.77142,
  63.06107, 62.74918, 62.758, 62.6357, 62.56111, 62.9577, 63.85057, 64.3729,
    64.43691, 64.24289, 64.01871, 63.44363, 61.34141, 61.50518, 60.52916,
    60.21236, 61.74081, 60.8713, 59.27539, 59.59624, 57.92038, 57.00873,
    58.89761, 59.5765, 59.4071, 59.17389, 59.21491, 59.17403, 58.36967,
    42.60637,
  64.63177, 63.50415, 63.2862, 63.08652, 63.00949, 63.37971, 63.68339,
    62.61168, 57.96788, 60.21488, 60.26173, 59.97043, 60.34615, 60.83939,
    61.19738, 61.16119, 60.758, 59.76812, 58.28347, 57.09685, 56.66977,
    57.04634, 58.41165, 59.4446, 59.37144, 59.51553, 59.51963, 58.92935,
    55.12167, 42.81525,
  68.35207, 66.45756, 65.0054, 64.2527, 63.87859, 63.50718, 62.37979,
    62.39123, 61.73856, 59.46414, 58.82952, 58.63441, 58.78951, 60.44463,
    61.87418, 61.62762, 62.42929, 62.49226, 62.08434, 61.09294, 60.24737,
    59.69608, 59.26297, 58.75932, 58.85545, 59.59989, 59.76625, 58.59959,
    42.83408, 43.27133,
  72.98155, 71.92587, 69.5955, 67.61523, 66.31812, 64.63928, 62.70108,
    62.83267, 62.63815, 62.37177, 60.95855, 58.85488, 57.4425, 56.36711,
    56.13158, 57.1772, 58.59603, 60.11895, 61.3637, 61.52051, 61.19734,
    60.25988, 59.28767, 58.51511, 58.59933, 58.84048, 58.74613, 47.96283,
    42.77446, 42.8261,
  75.36327, 75.33099, 76.06731, 73.50621, 71.34765, 67.65493, 65.23109,
    63.78938, 63.09043, 63.26703, 62.01944, 60.80118, 58.54626, 55.64188,
    53.64398, 53.54591, 53.18165, 53.32771, 54.38943, 56.3993, 59.52208,
    60.22385, 59.1591, 59.05796, 59.61047, 59.21526, 50.37972, 43.12376,
    43.60908, 42.90206,
  73.95448, 73.4724, 76.80067, 78.31705, 76.78798, 72.67569, 68.45029,
    64.85727, 63.24856, 63.22403, 62.53237, 61.75762, 61.40963, 61.14817,
    60.51088, 56.91838, 56.48779, 54.84548, 53.43582, 53.48791, 56.06351,
    57.17923, 56.29857, 58.74563, 59.01139, 58.58388, 43.35289, 47.2538,
    44.17899, 43.39137,
  65.66293, 67.39595, 69.21989, 71.94017, 74.16483, 74.0158, 68.15182,
    63.59355, 65.57044, 64.13811, 63.59233, 62.81599, 62.74157, 62.5589,
    61.7397, 60.14068, 60.19543, 60.22679, 60.05892, 56.72982, 57.40568,
    58.59178, 56.36366, 51.10136, 50.07, 51.05467, 43.55974, 45.13286,
    44.88366, 43.971,
  64.39025, 64.02464, 63.77632, 62.95932, 63.02863, 64.00578, 65.35869,
    65.91468, 64.05843, 64.33336, 64.19317, 63.35375, 63.0024, 62.85028,
    61.96644, 60.87926, 60.42553, 60.59216, 60.73652, 59.92355, 59.30455,
    55.77335, 48.62029, 45.45741, 43.133, 43.41012, 43.4557, 42.98053,
    43.26496, 43.39643,
  65.68259, 64.2906, 65.10736, 64.44915, 64.09682, 64.30329, 64.83614,
    64.78098, 64.10181, 63.59702, 63.14703, 62.65182, 62.67307, 62.3749,
    61.88283, 61.73008, 60.90015, 60.65865, 59.16642, 55.42274, 49.04416,
    49.35841, 46.95749, 43.83622, 44.61523, 44.20421, 43.63272, 43.17211,
    42.88083, 42.89448,
  60.67216, 62.38027, 62.70293, 63.1951, 63.49937, 64.59467, 64.98633,
    64.96315, 64.50074, 63.83847, 63.58827, 63.39575, 63.3324, 63.50315,
    62.56266, 61.72065, 61.52847, 56.86953, 52.45144, 50.22613, 48.17799,
    47.02377, 44.97705, 44.12349, 44.23691, 44.15706, 43.55952, 43.12722,
    42.95332, 42.98057,
  62.02969, 61.00755, 60.96744, 60.96471, 60.87414, 60.92781, 61.72043,
    63.65113, 64.59969, 64.20844, 63.87753, 64.40167, 65.14829, 64.97752,
    64.19823, 63.78581, 63.40766, 60.55909, 56.26068, 52.63557, 48.71519,
    47.76202, 45.74791, 44.53862, 44.55322, 44.2795, 43.49183, 42.93181,
    42.86394, 42.90245,
  68.77238, 65.16509, 62.42931, 61.46666, 61.30464, 60.68191, 60.56717,
    60.89393, 61.48683, 60.86092, 61.8757, 63.45584, 64.49474, 64.4325,
    64.25399, 64.91221, 65.7643, 66.01037, 64.93655, 59.83927, 52.95843,
    49.06045, 46.81453, 45.68611, 44.93797, 44.47719, 43.6855, 42.93892,
    42.80848, 42.87236,
  80.41652, 75.77869, 67.1088, 61.65603, 62.65475, 61.58833, 61.37335,
    61.15563, 60.25032, 59.96679, 59.763, 58.71013, 56.55995, 55.85603,
    55.82479, 58.00255, 62.29781, 65.85494, 66.10713, 65.2318, 60.12803,
    52.94776, 48.63392, 47.57772, 46.13268, 45.30874, 44.3922, 43.15015,
    42.79949, 42.85513,
  80.22498, 76.50841, 68.66557, 63.80186, 64.59475, 63.89024, 63.48041,
    63.0413, 62.85254, 62.76478, 62.3221, 60.87187, 59.81551, 56.54762,
    53.92509, 52.98958, 53.94873, 56.16114, 57.49581, 58.08433, 57.37191,
    54.48571, 50.56621, 48.95496, 47.31697, 45.9556, 44.81156, 43.38295,
    42.7172, 42.86979,
  79.8992, 77.19361, 69.96304, 65.86997, 66.88275, 66.33182, 66.21412,
    65.98572, 65.65477, 65.01563, 63.53975, 62.04156, 61.83588, 60.50746,
    58.36542, 57.23774, 56.32978, 55.93248, 55.41624, 53.90361, 53.05193,
    52.89952, 51.93334, 49.89198, 48.50953, 46.64597, 44.98389, 43.42536,
    42.71343, 42.85637,
  78.6167, 76.88542, 70.18473, 66.74961, 68.66949, 68.62548, 69.06054,
    69.38669, 69.90606, 69.61125, 68.08487, 66.30567, 64.99073, 63.53267,
    61.95817, 60.613, 59.30814, 58.17905, 57.01087, 54.73407, 52.03527,
    50.9303, 52.53513, 50.55358, 49.69917, 47.46706, 45.55011, 43.94933,
    42.9137, 42.84487,
  77.33298, 76.09034, 69.38196, 66.08579, 68.55344, 69.62776, 70.54756,
    71.18205, 72.71152, 73.49671, 73.36834, 73.28082, 72.44358, 71.12974,
    69.24573, 67.37805, 65.4727, 63.44683, 61.58028, 58.6631, 55.02088,
    52.71436, 52.83316, 51.33419, 51.22141, 49.10921, 46.5945, 44.87067,
    43.65865, 43.02688,
  76.3371, 73.90373, 67.73459, 65.01651, 66.82002, 67.63414, 69.23464,
    71.26482, 74.28612, 75.85284, 76.26224, 78.33445, 79.16858, 79.27888,
    77.93966, 76.42381, 73.53889, 70.65778, 67.78331, 64.54733, 61.37032,
    58.10322, 55.05253, 53.40159, 52.8787, 51.65082, 49.30545, 46.1014,
    44.73381, 43.66203,
  75.27174, 71.06863, 63.83356, 60.47348, 61.23877, 61.9972, 64.5845,
    68.12092, 72.28559, 72.61126, 73.01922, 75.15951, 78.01295, 78.62467,
    77.29155, 76.08405, 73.82745, 71.3072, 69.10484, 66.62132, 63.25338,
    60.0082, 56.49809, 54.18561, 53.7005, 52.40687, 50.68993, 47.30869,
    45.00928, 44.14278,
  74.43747, 69.65535, 63.37077, 59.11709, 58.88261, 58.54184, 60.83649,
    64.72609, 67.52079, 67.50932, 69.2484, 71.78022, 74.58303, 75.50672,
    73.85181, 72.739, 71.04558, 69.07297, 67.41658, 65.94357, 63.57915,
    60.85614, 57.29927, 54.9618, 54.66945, 53.19181, 51.66136, 48.43322,
    44.89825, 43.76737,
  71.6805, 67.30879, 61.72706, 57.83207, 57.713, 56.56693, 57.27508,
    58.84352, 60.3432, 60.57912, 62.53883, 65.15281, 68.29402, 69.52357,
    68.82888, 68.03776, 66.515, 65.09705, 64.34988, 63.31546, 62.00975,
    59.49692, 56.58723, 54.79295, 54.64553, 53.72511, 52.83445, 50.21314,
    46.16362, 43.68626,
  64.33417, 62.41979, 58.38141, 55.86726, 56.98123, 56.49113, 55.37688,
    54.58825, 54.01557, 53.95335, 54.60882, 56.08448, 58.45914, 60.10758,
    60.00227, 59.39402, 58.58402, 57.64929, 57.37662, 58.15066, 57.26326,
    55.60498, 53.06, 51.63641, 51.80066, 51.29303, 50.36051, 49.38477,
    47.50182, 44.48699,
  49.95969, 50.84056, 51.58455, 52.20591, 53.29297, 54.76782, 52.86848,
    49.74081, 48.86804, 49.09472, 48.65921, 48.38706, 48.49148, 48.98115,
    48.97495, 48.89968, 48.27546, 47.87676, 47.73677, 47.76043, 48.37584,
    49.00947, 49.03088, 48.36407, 48.41799, 48.16214, 47.38253, 45.85468,
    44.98946, 44.27193,
  46.40696, 46.7948, 47.30857, 47.27581, 47.94796, 49.51307, 49.7107,
    47.32093, 46.19782, 46.626, 46.74845, 46.8123, 46.55748, 46.23647,
    45.99088, 45.72437, 44.98965, 44.16471, 44.03689, 44.10033, 44.01473,
    44.58799, 45.44878, 45.86474, 45.75418, 45.82253, 45.36877, 44.42075,
    43.67767, 43.07941,
  56.85157, 56.68154, 56.30941, 55.93447, 55.35276, 54.88975, 54.51488,
    54.34522, 54.45432, 54.95424, 56.02703, 57.02877, 57.24504, 58.12236,
    58.89566, 58.9033, 58.80556, 58.47364, 57.50339, 56.30251, 54.62965,
    52.48754, 51.38577, 51.30249, 50.74004, 47.8649, 45.73059, 47.19188,
    43.56186, 41.95446,
  59.99921, 60.10996, 59.70982, 59.51357, 58.88352, 58.22599, 57.66591,
    57.07719, 56.47975, 56.06161, 56.2472, 57.10715, 58.20832, 59.04008,
    59.28923, 59.34647, 59.35223, 59.42535, 59.50567, 59.57172, 59.51065,
    59.35369, 59.18067, 59.38024, 59.44636, 57.23448, 44.04801, 45.65917,
    43.4731, 42.23362,
  60.42908, 60.3144, 60.26042, 60.1559, 59.95119, 59.81453, 59.71442,
    59.65398, 59.601, 59.42562, 59.24916, 58.45648, 57.82678, 57.6252,
    57.82447, 57.91748, 59.19873, 59.40216, 59.71091, 60.02831, 60.52169,
    60.92915, 60.97747, 60.88173, 60.27003, 58.75892, 56.43103, 46.56742,
    42.83416, 42.36114,
  60.65554, 60.6376, 60.60572, 60.51811, 60.36381, 60.21614, 60.13578,
    60.03741, 59.94333, 59.74365, 59.77538, 60.13531, 60.22737, 59.96693,
    59.89198, 59.82484, 59.43681, 59.2272, 59.54333, 60.04922, 60.50084,
    60.44843, 60.51342, 60.96469, 60.4071, 59.40904, 58.61966, 57.93425,
    48.82127, 43.17965,
  60.75097, 60.77641, 60.7952, 60.70526, 60.46509, 60.48766, 60.55734,
    60.27351, 59.99852, 59.68296, 59.84651, 60.63591, 61.18085, 61.06716,
    61.1094, 61.2661, 60.70868, 59.75481, 59.69535, 60.12706, 59.96582,
    57.70196, 58.41396, 60.01748, 60.1772, 59.70422, 59.45791, 59.93523,
    59.55563, 51.59418,
  60.56542, 60.7597, 60.87505, 60.82689, 60.58513, 60.88491, 61.50779,
    61.37579, 60.87579, 60.44936, 60.43115, 61.12571, 61.83895, 61.72235,
    62.17706, 62.70455, 61.99583, 60.77958, 59.90517, 59.86431, 59.52121,
    54.01783, 58.03627, 59.61146, 59.6572, 59.74121, 60.02953, 60.60494,
    59.56881, 45.74076,
  60.34201, 60.44941, 60.63859, 60.66531, 60.55775, 61.05599, 62.02121,
    62.27454, 62.03946, 61.65494, 61.27694, 60.61129, 58.23785, 58.89813,
    59.28107, 60.39862, 60.29633, 59.40287, 58.83002, 58.99068, 58.13963,
    57.00021, 58.8344, 59.76726, 59.6091, 59.40919, 59.93895, 60.04316,
    58.31168, 41.08846,
  60.48697, 60.31869, 60.44747, 60.39169, 60.41217, 60.92733, 61.38682,
    60.54346, 58.71619, 60.24168, 60.18885, 59.51799, 59.10239, 59.05806,
    59.11729, 59.15166, 59.19816, 58.61235, 57.33666, 56.79553, 57.3345,
    58.86362, 59.66326, 59.81762, 59.56197, 59.67899, 60.092, 59.50244,
    52.38095, 41.29814,
  61.95626, 61.29409, 60.84826, 60.58009, 60.30791, 60.12461, 57.90179,
    56.39066, 57.37246, 57.73603, 58.77972, 59.75686, 60.23375, 60.751,
    61.13662, 60.88983, 61.12859, 61.38251, 61.17704, 60.29533, 59.67419,
    59.73466, 59.76383, 59.44672, 59.44717, 60.02763, 59.80663, 58.50705,
    41.54609, 41.85231,
  64.92432, 64.18569, 63.11129, 62.32618, 61.71914, 60.48455, 57.74674,
    59.47472, 58.14319, 56.81477, 55.93159, 56.6911, 56.80574, 56.8529,
    57.35103, 59.82333, 60.59172, 60.9831, 61.14823, 61.0786, 60.93334,
    60.21491, 59.33668, 58.62239, 59.24102, 59.87716, 58.94243, 46.88776,
    41.29124, 41.24506,
  69.03678, 67.8792, 68.44086, 66.2628, 65.4328, 62.72638, 61.0888, 60.07551,
    59.93904, 60.23794, 57.5197, 52.41608, 51.62633, 50.8753, 50.61451,
    51.43335, 52.40409, 53.65595, 55.59372, 58.95622, 60.76744, 60.41139,
    59.20673, 58.87985, 59.29537, 58.90553, 48.95205, 41.59953, 42.19945,
    41.3397,
  73.39635, 71.9353, 73.61412, 73.73901, 71.06371, 67.37057, 64.12288,
    61.07943, 59.36777, 59.84747, 59.3288, 58.61409, 58.62377, 58.52034,
    55.77069, 53.01868, 53.00122, 52.429, 52.29349, 53.71836, 58.14809,
    60.12028, 59.1154, 59.33156, 59.41888, 58.21278, 42.13087, 45.71843,
    42.77499, 41.85134,
  65.85178, 67.65495, 69.36395, 71.08306, 71.85613, 69.82871, 63.20637,
    60.02104, 61.63599, 60.46944, 60.1673, 59.65893, 59.83617, 60.02068,
    59.67553, 57.60809, 58.72333, 59.06815, 58.08596, 55.78833, 57.68605,
    59.20044, 56.84104, 52.22807, 51.81073, 49.66053, 42.53506, 44.07386,
    43.64971, 42.51845,
  61.00188, 60.98053, 61.00652, 60.09193, 60.13474, 60.83388, 61.86753,
    61.95469, 60.21924, 60.61906, 60.73312, 60.00353, 59.97905, 60.25221,
    59.63261, 58.9252, 58.89569, 59.47343, 59.98298, 59.57574, 59.49847,
    57.70047, 50.77693, 44.87827, 41.89547, 42.30823, 41.99755, 41.66367,
    41.99454, 41.98389,
  63.23544, 62.70624, 62.34892, 61.36576, 60.71476, 60.6823, 61.38077,
    61.21377, 59.74693, 59.59808, 59.36856, 59.24602, 59.60409, 59.56768,
    59.47376, 59.47805, 58.87614, 59.23563, 59.63824, 58.47315, 52.12038,
    49.7646, 45.05676, 42.91199, 43.4221, 42.91983, 42.26342, 41.77298,
    41.48322, 41.42842,
  58.69957, 61.31941, 62.28555, 62.12921, 61.95452, 62.33646, 62.55059,
    62.22918, 61.46574, 60.42198, 59.61013, 58.66097, 58.57242, 59.99096,
    58.12707, 57.11078, 57.89547, 53.76423, 50.799, 48.5994, 46.16332,
    45.70317, 43.68283, 42.84489, 43.11579, 42.97179, 42.21174, 41.8173,
    41.57952, 41.47382,
  55.70721, 55.45752, 56.23201, 57.30551, 58.49223, 59.71474, 61.49637,
    62.45231, 62.40983, 61.85827, 61.30344, 61.57421, 62.22513, 61.90937,
    60.78777, 59.88179, 57.44133, 55.36403, 52.99826, 50.30136, 46.39817,
    46.11946, 44.1875, 43.1872, 43.24354, 43.05184, 42.08441, 41.448,
    41.40276, 41.41048,
  60.12846, 57.38935, 55.13049, 54.78729, 55.22511, 55.95393, 57.21537,
    59.04091, 60.75718, 61.43581, 62.22643, 62.70181, 62.95584, 62.89492,
    62.52421, 62.76802, 63.30162, 63.58198, 61.39838, 56.2971, 49.66227,
    46.86085, 45.18495, 44.24755, 43.4796, 42.89524, 42.15846, 41.37637,
    41.30518, 41.31161,
  75.07538, 67.55986, 58.66488, 53.43952, 54.31153, 53.67456, 54.05717,
    54.58784, 54.60183, 55.41858, 56.84218, 56.90636, 55.68829, 56.53448,
    57.25066, 59.69734, 63.67044, 65.2253, 65.3055, 64.01132, 57.28637,
    50.55498, 46.95494, 45.94679, 44.50234, 43.50507, 42.59029, 41.55409,
    41.29181, 41.34649,
  75.98817, 69.81347, 61.20615, 55.92696, 56.21482, 55.44661, 55.29234,
    55.24901, 55.50526, 56.16117, 56.06875, 54.5765, 54.3748, 52.47436,
    50.93282, 50.9321, 53.01321, 56.41233, 57.97702, 58.06891, 56.16717,
    52.61668, 48.96897, 47.33812, 45.71213, 44.07954, 42.91327, 41.721,
    41.23568, 41.3485,
  77.2246, 73.18424, 64.70197, 59.92852, 59.95734, 58.86997, 58.39802,
    58.07329, 57.94941, 57.54777, 55.96646, 54.64311, 55.5409, 54.87825,
    53.41112, 52.92238, 53.19916, 53.91278, 54.3373, 53.20989, 52.46777,
    52.09718, 50.64256, 48.71418, 46.7791, 44.64029, 43.0342, 41.79276,
    41.24183, 41.33368,
  77.23049, 75.40803, 68.28291, 64.60629, 65.33165, 64.32822, 63.89519,
    63.28172, 63.29255, 62.31767, 59.88991, 58.21704, 57.68579, 56.81328,
    55.71783, 55.01929, 54.45663, 54.45766, 54.45456, 53.86221, 52.97379,
    51.48981, 50.67429, 49.80401, 48.17718, 45.55996, 43.56103, 42.29601,
    41.39283, 41.31323,
  76.43794, 75.1861, 69.2992, 66.49073, 68.52942, 68.9054, 68.85087,
    68.41228, 69.16173, 68.68163, 67.05128, 66.98978, 66.06225, 64.43664,
    62.49029, 61.08047, 59.52101, 57.79584, 56.48305, 55.14353, 53.75318,
    51.97434, 50.44626, 50.12123, 50.11438, 47.70913, 44.85069, 43.24553,
    42.13751, 41.44355,
  75.20418, 73.33144, 68.55393, 66.21133, 67.35289, 67.51656, 68.6439,
    70.39857, 73.22308, 74.08166, 73.15344, 74.979, 75.68265, 75.13998,
    73.2168, 71.23809, 68.61784, 65.62397, 62.6487, 59.95128, 57.47866,
    55.07498, 52.72853, 51.52452, 51.53577, 50.78077, 48.05496, 44.72406,
    43.36023, 42.14604,
  74.20226, 70.71815, 64.2691, 61.28931, 61.58148, 61.8864, 64.4489,
    68.74883, 73.32651, 72.71498, 71.35095, 73.16765, 75.04784, 75.31877,
    73.7377, 72.36935, 69.79432, 67.35742, 65.46173, 63.29644, 60.3855,
    57.4831, 54.22977, 52.10823, 52.03312, 51.41427, 49.99222, 46.38635,
    44.01555, 42.76544,
  72.29142, 69.12615, 63.68451, 59.75984, 58.89245, 58.49008, 61.47291,
    66.4177, 69.75624, 68.70236, 69.6107, 71.42887, 73.35576, 73.46378,
    71.8865, 70.62592, 68.6216, 66.47169, 65.35997, 64.29969, 62.2407,
    59.58958, 56.29115, 53.93464, 53.53825, 52.32735, 50.90796, 47.54181,
    43.58338, 42.29206,
  70.14993, 66.56796, 61.51179, 57.9931, 57.38666, 56.07867, 57.71539,
    60.23711, 62.09402, 62.14222, 63.91505, 66.37876, 68.7298, 69.46042,
    68.40813, 67.51819, 65.75591, 64.11297, 63.72864, 63.19073, 61.40398,
    59.52278, 57.12968, 55.38061, 55.03242, 54.30304, 53.4986, 50.6136,
    44.99181, 42.02604,
  64.34125, 62.04274, 58.86326, 56.83428, 57.74468, 56.94709, 55.89154,
    55.59309, 54.67146, 54.99452, 55.75279, 57.48388, 59.79167, 60.90467,
    60.56042, 60.22343, 59.01128, 58.22773, 58.47523, 58.94843, 57.57083,
    55.07961, 52.69559, 51.3215, 51.62504, 51.37787, 50.75212, 50.10573,
    47.58796, 43.18649,
  50.79725, 51.6074, 52.2212, 52.8815, 54.57513, 56.26818, 53.91355,
    50.03059, 49.05576, 49.41772, 49.07188, 48.80154, 48.87216, 49.2999,
    49.35921, 49.31782, 48.79099, 48.28064, 48.08772, 48.056, 48.15076,
    48.46571, 48.08447, 47.2187, 47.40517, 47.35128, 46.6128, 45.07101,
    44.3518, 43.20441,
  46.40147, 46.87197, 47.22632, 47.10229, 48.06575, 50.21328, 50.54169,
    47.2085, 45.71395, 46.58968, 47.05337, 47.19778, 46.88348, 46.43209,
    45.96569, 45.57379, 44.48212, 43.31882, 43.21852, 43.25868, 43.0864,
    43.64784, 44.40578, 44.73145, 44.64012, 44.82847, 44.40657, 43.25307,
    42.30242, 41.54708,
  51.47485, 51.63708, 51.86231, 52.34314, 52.70854, 53.16056, 53.72869,
    54.31191, 54.92248, 55.76377, 56.91711, 56.74671, 54.49146, 54.17812,
    53.91096, 53.12349, 52.85149, 53.07047, 53.12567, 53.45945, 53.06615,
    51.38758, 51.48363, 53.01851, 53.80735, 52.11292, 52.72073, 53.84003,
    45.12276, 42.19562,
  55.32627, 55.37001, 54.83141, 55.3186, 55.12864, 55.23354, 55.95666,
    56.76924, 57.7206, 58.87027, 59.67792, 60.06639, 60.29387, 60.09465,
    59.96804, 60.10682, 60.11355, 60.40015, 60.68411, 60.88107, 60.8091,
    60.57783, 60.52101, 61.01463, 61.20493, 58.48803, 49.11192, 51.62067,
    45.25195, 42.94014,
  57.86719, 58.24648, 58.30164, 58.23253, 58.00588, 57.8733, 57.85899,
    58.04444, 58.23523, 58.53069, 59.19996, 60.0214, 60.37169, 60.72789,
    60.92422, 60.68734, 60.76596, 61.10174, 61.4528, 61.80571, 62.26545,
    62.65594, 62.69707, 62.74251, 62.27282, 60.63341, 58.64318, 50.93861,
    44.63392, 43.39633,
  59.51562, 59.58069, 59.79964, 59.97273, 60.02406, 60.15304, 60.31159,
    60.41006, 60.39862, 60.23328, 60.30057, 60.72898, 60.93887, 60.84435,
    61.31044, 61.54345, 61.06806, 60.73097, 61.27971, 62.01093, 62.70766,
    62.82902, 63.10776, 63.76816, 63.18829, 61.81224, 60.32499, 59.22452,
    48.67272, 43.31347,
  59.98458, 59.9251, 60.07962, 60.14393, 60.05655, 60.17643, 60.55257,
    60.64185, 60.63326, 60.51219, 60.57154, 61.35649, 62.01867, 62.09368,
    62.28372, 62.6284, 62.12798, 60.9847, 61.07766, 61.863, 61.94908,
    61.5131, 62.03953, 62.97878, 63.34254, 62.35989, 60.97432, 61.0442,
    60.75722, 51.47517,
  60.13007, 60.45435, 60.77267, 60.89678, 60.5316, 60.68601, 61.41378,
    61.37788, 61.01058, 60.87669, 61.15081, 62.17659, 63.19812, 63.19977,
    63.86216, 64.4838, 63.83592, 62.50901, 61.34792, 61.68368, 61.48089,
    58.9889, 61.71321, 62.36742, 62.69834, 62.26667, 61.58818, 62.10723,
    61.02745, 46.61797,
  60.10496, 60.57802, 61.00465, 61.22796, 61.07116, 61.48729, 62.41048,
    62.57596, 62.21655, 61.91466, 61.79596, 61.49161, 61.06547, 61.60669,
    62.2257, 62.76417, 62.7428, 61.73618, 60.80083, 61.2439, 61.36169,
    61.60228, 62.11726, 62.76825, 62.54857, 61.57541, 61.69965, 61.6421,
    59.96115, 41.19025,
  60.34163, 60.69995, 61.2674, 61.70612, 61.76208, 62.41615, 63.12119,
    62.4467, 61.90057, 62.09206, 62.08036, 62.14934, 62.30568, 62.56599,
    62.86605, 63.28648, 63.498, 63.14779, 62.2611, 61.86579, 61.96377,
    62.52086, 63.21949, 63.40562, 62.50949, 62.08299, 62.37951, 61.60387,
    56.14816, 41.81874,
  62.02569, 62.10601, 62.10709, 62.04872, 61.71826, 61.81503, 61.7565,
    62.59901, 63.35748, 63.7178, 63.92347, 64.04819, 64.40137, 65.6711,
    66.3186, 65.04441, 65.29787, 65.79615, 65.48164, 63.96705, 63.04182,
    63.72533, 64.46735, 63.78621, 62.65867, 63.19825, 62.31274, 60.58388,
    43.34666, 42.29471,
  64.34648, 64.93727, 64.17414, 64.22632, 63.46807, 62.01909, 60.81487,
    61.80238, 62.27348, 63.09439, 63.60613, 63.87478, 63.65059, 63.49409,
    63.31544, 64.46131, 65.05072, 65.34613, 65.39667, 65.36527, 65.23553,
    64.06228, 62.60542, 61.05288, 61.55484, 62.24009, 60.97551, 49.86772,
    41.66778, 40.75317,
  65.1224, 64.79377, 65.90939, 64.74886, 65.45624, 63.72461, 62.6474,
    62.30448, 63.01597, 63.83265, 62.30113, 57.33984, 55.41447, 55.77723,
    56.11448, 57.89205, 59.90208, 61.32617, 62.03166, 62.96124, 64.51579,
    63.49939, 60.9627, 60.15382, 60.50726, 60.12721, 49.95301, 42.1807,
    42.48018, 40.9086,
  70.01659, 67.86327, 69.81705, 70.58098, 68.58121, 66.35163, 64.3619,
    62.00016, 60.50662, 61.13653, 60.87346, 59.9855, 60.71043, 61.18984,
    57.97116, 57.88753, 57.35559, 57.47219, 57.89599, 60.8793, 63.14021,
    62.97381, 60.71257, 61.11327, 60.9341, 59.44186, 42.56549, 46.36293,
    43.48465, 41.86197,
  68.53027, 69.87991, 71.4858, 72.7997, 72.73869, 70.62976, 64.47324,
    61.23451, 62.98963, 61.89985, 62.22125, 62.01057, 62.88113, 63.18723,
    61.60326, 60.59951, 60.84573, 61.15215, 61.33894, 62.06157, 62.73014,
    62.14388, 60.46192, 56.22562, 55.11485, 51.29863, 43.65379, 45.17026,
    44.83352, 42.86723,
  61.48815, 62.11258, 62.61463, 62.1232, 62.17574, 62.89758, 63.96896,
    64.21428, 62.75776, 63.93007, 64.85017, 64.29524, 65.03604, 64.92966,
    63.42289, 61.71025, 61.09151, 61.74437, 62.33405, 62.14624, 61.71034,
    60.45227, 53.76263, 47.35509, 44.14163, 43.8143, 42.59854, 42.05041,
    42.43731, 42.13689,
  62.75122, 63.2493, 62.8077, 62.3443, 62.38839, 64.01568, 65.92418,
    64.54217, 62.98548, 62.67019, 62.25019, 61.93897, 62.32867, 63.22332,
    62.87542, 61.613, 61.33199, 62.00803, 62.9665, 62.48464, 55.81572,
    53.08242, 47.2431, 45.2078, 45.29899, 44.26896, 42.99852, 42.11692,
    41.51252, 41.23248,
  62.64563, 63.38955, 63.62045, 63.33926, 63.10811, 63.79661, 64.62095,
    64.23666, 63.01431, 61.97882, 61.81314, 61.22257, 60.99726, 61.89588,
    61.40166, 60.9356, 61.36478, 61.64485, 60.90007, 56.48234, 49.74166,
    49.69308, 45.86398, 44.67538, 44.83239, 44.25949, 42.77195, 42.2491,
    41.73479, 41.30367,
  61.2836, 61.50078, 61.81645, 62.26377, 62.71652, 62.9204, 63.58833,
    64.59418, 64.56584, 63.77569, 62.73331, 63.34212, 64.62929, 63.78743,
    62.2351, 61.76976, 61.68844, 61.67037, 61.32701, 57.49723, 49.42581,
    49.89515, 46.69104, 44.89152, 44.53961, 44.20826, 42.44012, 41.34773,
    41.30927, 41.18806,
  58.85064, 58.54134, 57.99352, 59.81781, 61.6944, 62.19885, 62.90548,
    63.86588, 64.62136, 64.54129, 65.30595, 66.07585, 66.05243, 66.06737,
    65.15479, 64.83892, 64.84833, 65.31366, 65.05981, 62.94558, 51.70037,
    49.5129, 47.20567, 46.00146, 44.11625, 43.1226, 42.44902, 41.11049,
    41.06579, 40.96313,
  69.12885, 63.68063, 56.76997, 53.53391, 55.62019, 56.55422, 58.6022,
    60.88307, 62.26664, 63.25931, 64.07111, 64.02641, 63.43352, 63.93879,
    64.11059, 65.17847, 67.52819, 69.65386, 69.43148, 67.36678, 61.81183,
    53.31954, 48.87189, 47.04716, 44.67344, 43.21741, 42.43232, 41.38447,
    41.04882, 40.98101,
  68.81585, 63.7252, 56.96286, 52.8833, 54.03045, 54.59723, 55.80938,
    57.18874, 59.33876, 62.6566, 62.75613, 58.73281, 59.28628, 58.60574,
    57.51949, 57.62254, 61.14519, 64.93865, 66.01105, 65.84299, 64.53861,
    58.39755, 52.07434, 48.97152, 46.53729, 43.96433, 42.66188, 41.52767,
    41.00931, 40.99156,
  70.78571, 65.94653, 58.59382, 54.56476, 54.68506, 54.61969, 55.28753,
    56.3528, 58.20153, 59.77553, 57.401, 54.47541, 57.24535, 57.2424,
    56.11975, 55.50316, 56.42708, 57.88874, 59.67756, 59.71946, 59.7217,
    59.87877, 56.8723, 52.61869, 48.60168, 45.03574, 42.77774, 41.5565,
    40.97948, 41.0159,
  73.14684, 70.87601, 64.34679, 61.05241, 61.22192, 59.77387, 59.90421,
    60.01009, 61.72516, 61.53248, 57.21902, 55.22801, 56.52843, 56.32389,
    55.60688, 55.57323, 55.27145, 55.527, 56.56438, 57.11391, 57.66402,
    57.35424, 57.50188, 56.71514, 52.36374, 46.49634, 43.39325, 42.31776,
    41.21667, 40.97154,
  74.58745, 73.44158, 69.16311, 67.2626, 68.03252, 67.99801, 67.80705,
    67.24279, 67.95002, 66.36462, 62.33077, 63.1434, 63.47984, 62.99168,
    61.32211, 60.73572, 59.69047, 57.29002, 56.31744, 55.9516, 55.65794,
    54.92733, 54.25676, 55.28849, 55.76392, 50.70712, 45.59276, 44.01443,
    42.45713, 41.14544,
  74.99007, 73.69045, 70.34042, 68.81866, 69.18414, 69.00413, 69.60511,
    70.73679, 72.9063, 73.03874, 70.85342, 73.295, 74.36187, 74.28985,
    73.15291, 71.84765, 69.40381, 65.90794, 62.14962, 59.89893, 58.27527,
    56.7237, 55.18256, 54.82266, 55.91691, 55.98221, 51.48112, 46.29341,
    44.45613, 42.20319,
  74.90021, 72.43331, 68.43932, 66.57551, 66.73517, 66.63, 68.33714,
    71.16959, 74.11923, 73.51419, 71.32024, 73.64773, 74.88578, 75.19754,
    74.39577, 73.81946, 72.71667, 70.57382, 68.27682, 65.75729, 62.85201,
    59.90659, 56.94638, 55.10918, 55.52958, 56.43876, 55.45904, 50.09445,
    46.33804, 43.837,
  74.45675, 72.22665, 68.62085, 66.30925, 65.95474, 65.01859, 67.9746,
    71.31853, 73.31802, 72.51547, 72.88761, 73.74658, 74.87207, 74.82964,
    73.8754, 73.48358, 72.83691, 71.83768, 71.05923, 70.06223, 68.27363,
    65.9054, 62.14961, 59.20275, 58.7801, 57.8301, 56.99922, 52.0063,
    44.93598, 42.84712,
  72.42963, 70.28594, 67.19612, 65.25602, 65.23476, 63.28601, 66.0789,
    68.73212, 68.88625, 67.87181, 70.52555, 72.43221, 73.64276, 73.77316,
    72.57236, 71.6303, 70.91669, 70.59072, 70.4417, 69.82281, 69.12826,
    68.63908, 67.36587, 65.78795, 65.12787, 64.16244, 63.84775, 59.57571,
    48.09805, 41.79618,
  68.49667, 67.18038, 65.19146, 64.15151, 64.88653, 64.89754, 65.20411,
    63.90178, 60.558, 61.37941, 62.81976, 64.93023, 67.01325, 67.8727,
    67.91576, 67.26733, 65.45615, 64.96492, 65.70462, 66.2274, 63.94889,
    60.8189, 58.41073, 57.93755, 58.95136, 59.23539, 59.158, 60.21244,
    55.79165, 44.81792,
  59.26281, 60.07662, 60.8279, 61.26574, 62.53384, 63.93507, 63.45849,
    57.8943, 55.37496, 56.30425, 55.95057, 56.10987, 56.77365, 57.44203,
    57.91637, 57.72124, 56.51943, 55.61496, 54.37544, 52.6223, 51.90834,
    51.44566, 50.13997, 49.09986, 49.99722, 50.83078, 50.34283, 48.38392,
    47.8609, 45.42125,
  52.78682, 53.29635, 53.47328, 53.15999, 55.37881, 60.56373, 62.23272,
    54.34639, 50.67794, 52.95107, 54.50728, 55.93681, 55.87886, 54.88459,
    53.44245, 52.37464, 49.2001, 46.09316, 45.74482, 45.33904, 44.31429,
    44.88298, 45.44659, 45.62034, 45.91043, 46.70021, 46.61173, 44.55879,
    42.53084, 41.01141,
  46.07499, 46.18618, 46.35398, 46.6186, 46.60413, 46.73, 47.06223, 47.57449,
    48.23267, 49.17689, 51.28194, 51.1245, 47.48465, 47.91222, 48.24231,
    47.64949, 47.83866, 48.7125, 49.83355, 51.71405, 52.38731, 50.89099,
    51.51483, 54.10615, 56.09644, 55.91116, 60.77901, 62.37293, 47.96862,
    44.30415,
  49.67949, 50.08425, 49.38514, 50.2272, 49.65832, 49.32577, 49.8051,
    50.37455, 50.98824, 51.7596, 53.1866, 55.03435, 56.00176, 53.74776,
    52.17986, 52.90673, 51.9015, 53.0114, 54.83357, 56.27882, 55.87476,
    55.04392, 55.56069, 59.2671, 62.5168, 58.31049, 56.03437, 60.2788,
    48.99694, 45.53296,
  49.10698, 49.80248, 50.68583, 51.33949, 51.85644, 52.31346, 52.36913,
    52.67999, 53.12572, 53.69868, 54.48963, 55.87609, 57.34699, 59.22436,
    60.12248, 57.86166, 58.07726, 59.58739, 60.58849, 62.3872, 62.73603,
    62.94493, 63.11063, 63.62024, 63.54665, 62.30616, 62.07898, 58.62111,
    48.66226, 46.70403,
  52.24242, 53.00682, 54.45657, 55.8391, 57.37452, 58.93081, 58.6801,
    57.96377, 58.26918, 58.97777, 59.18822, 59.93707, 59.75093, 58.84375,
    62.07828, 63.57814, 61.30704, 58.48337, 61.17887, 62.89027, 63.31142,
    63.52105, 64.07021, 65.11491, 65.35247, 64.19899, 62.40975, 58.56982,
    50.00859, 45.16983,
  54.34849, 54.12413, 56.3032, 57.72919, 58.59742, 58.94043, 58.98166,
    58.89331, 60.12863, 61.08836, 61.52179, 62.5932, 63.15096, 63.38908,
    63.6257, 64.20193, 63.71867, 61.19808, 62.28151, 62.92922, 62.98629,
    60.75452, 62.58952, 64.66451, 65.73956, 64.57176, 62.00768, 61.85207,
    61.90644, 50.71496,
  56.07877, 58.35867, 61.75361, 62.2888, 61.9848, 61.92162, 62.60601,
    62.61275, 62.1367, 62.03308, 62.33128, 63.18997, 64.03392, 63.97048,
    64.64322, 65.73113, 65.57959, 64.00126, 62.26188, 62.71223, 62.61256,
    58.15202, 61.98241, 64.06924, 65.07198, 64.26556, 62.40536, 62.91507,
    62.41346, 49.16422,
  58.53101, 61.10221, 61.80245, 62.20966, 61.99044, 62.13619, 62.64631,
    62.64156, 62.16935, 62.13906, 62.30838, 62.44236, 62.46508, 63.16532,
    63.94206, 64.73386, 65.24638, 63.9689, 62.17461, 62.76326, 61.72062,
    61.10145, 63.70519, 64.96319, 64.91174, 63.18096, 62.81551, 62.7853,
    61.95205, 44.66835,
  59.00346, 61.14722, 61.89363, 62.40466, 62.1793, 62.54034, 63.23658,
    62.71465, 60.2371, 61.92047, 61.85229, 61.79192, 62.18312, 63.9393,
    64.75902, 65.56088, 66.33804, 66.02566, 64.52161, 64.00963, 63.80245,
    64.35944, 65.42882, 65.92532, 64.73579, 63.70435, 64.087, 63.62297,
    60.46069, 45.14747,
  62.95433, 63.18054, 63.65268, 63.53377, 62.727, 63.08329, 63.5252,
    64.21869, 65.11794, 65.82922, 66.35101, 66.74707, 67.42747, 70.15151,
    71.73107, 69.32275, 69.89947, 70.74646, 70.16608, 68.00448, 66.64601,
    67.7974, 69.44239, 68.33622, 65.69723, 66.28889, 65.12633, 63.22748,
    49.10302, 44.60308,
  67.99794, 69.44181, 68.94719, 69.43717, 67.76733, 65.93277, 64.73605,
    65.71274, 66.32792, 68.15148, 69.77512, 70.97726, 70.45838, 68.96986,
    67.50898, 69.00362, 69.98161, 70.18331, 70.04681, 71.03082, 71.59714,
    69.55548, 67.69321, 65.13794, 64.5452, 64.57916, 63.46222, 53.20485,
    44.4011, 42.13081,
  66.10181, 65.61536, 67.08849, 66.93736, 67.93557, 67.23161, 66.55794,
    66.58331, 67.56875, 68.07861, 66.2841, 61.90228, 60.39849, 60.69993,
    61.79697, 63.34342, 64.23387, 64.91068, 65.88411, 66.88955, 68.41465,
    67.52943, 63.17143, 60.68747, 61.72522, 61.61891, 51.35059, 44.55891,
    44.12115, 42.25684,
  70.52222, 68.03354, 71.15604, 71.81033, 69.94047, 68.15665, 66.77116,
    64.6506, 62.65775, 62.30606, 59.9179, 57.96377, 60.6191, 62.34534,
    61.82449, 61.63108, 61.48993, 63.41734, 64.55051, 65.75964, 66.91767,
    66.37811, 61.72198, 62.69512, 62.23121, 56.21385, 45.15014, 46.97706,
    45.43463, 43.35324,
  73.98593, 75.58944, 77.2818, 77.25969, 76.09217, 72.77648, 65.77591,
    62.93787, 64.17596, 62.24062, 62.61377, 62.22644, 63.18432, 64.10003,
    63.75293, 63.08969, 63.58857, 64.29275, 66.12278, 68.9506, 68.09975,
    64.72984, 61.49456, 58.90931, 58.01812, 52.23885, 46.10025, 46.91263,
    46.90495, 44.35841,
  66.13069, 66.79304, 67.21236, 66.26868, 65.89824, 66.60857, 67.9958,
    68.10585, 65.25627, 65.18896, 65.51579, 63.94509, 65.18292, 65.98546,
    64.52042, 63.42743, 63.34139, 63.76197, 64.5875, 65.03344, 64.22406,
    61.76406, 57.4588, 51.4543, 48.42684, 47.40516, 45.04023, 44.23113,
    44.67847, 43.72307,
  63.17289, 64.02012, 64.54648, 64.58739, 64.41595, 65.23741, 67.98573,
    68.4104, 66.02846, 65.58187, 64.76945, 64.39894, 65.2846, 65.60763,
    64.86318, 64.28251, 63.89682, 64.76595, 66.34612, 65.98267, 57.61771,
    56.31093, 51.22836, 49.79978, 49.0807, 47.33047, 45.50315, 44.13113,
    43.33018, 42.72884,
  64.45354, 65.49709, 66.44753, 66.15835, 65.27122, 66.18684, 67.87363,
    67.30964, 66.09106, 65.05736, 65.28676, 64.20126, 63.58626, 65.06363,
    64.48257, 64.09325, 64.61723, 64.86388, 65.74689, 64.91613, 52.45945,
    53.18568, 49.42204, 48.43221, 48.56014, 47.3845, 45.11668, 44.38896,
    43.47871, 42.76855,
  62.87738, 62.56242, 63.12694, 63.51145, 63.86872, 64.20945, 65.2665,
    66.62634, 66.65653, 66.01518, 64.59345, 65.80877, 68.36554, 66.83498,
    64.8251, 64.42448, 64.26856, 64.56189, 65.74741, 64.9889, 51.56084,
    53.64123, 50.3837, 48.51941, 47.93428, 47.50391, 44.6889, 43.08858,
    43.01904, 42.66588,
  61.3357, 62.40377, 62.3886, 62.92754, 63.42894, 64.04232, 64.36621,
    64.98972, 65.80062, 65.45372, 67.05837, 69.64258, 69.62439, 68.08698,
    67.33843, 66.253, 65.0829, 65.6954, 67.05383, 64.99254, 52.81798,
    51.53416, 49.76678, 48.94152, 46.47192, 45.27053, 44.56343, 42.54399,
    42.47351, 42.29016,
  66.70686, 63.86802, 59.50657, 57.76288, 59.48026, 60.30038, 62.23608,
    63.68551, 63.83226, 64.6107, 66.28069, 66.36039, 64.68768, 65.10918,
    65.42483, 66.67908, 69.33865, 72.16289, 72.91071, 69.52445, 63.55068,
    54.16724, 50.47545, 48.82229, 45.98185, 44.4488, 43.88365, 42.78058,
    42.46473, 42.29814,
  64.71996, 62.56146, 59.2177, 56.45284, 57.73286, 58.57504, 59.39348,
    60.63986, 63.61063, 65.51125, 66.21931, 64.4436, 64.53751, 64.37114,
    63.85862, 64.81104, 66.97063, 69.03841, 68.60411, 67.94715, 66.27073,
    60.64354, 53.398, 50.62804, 48.15245, 45.13596, 43.97761, 42.92241,
    42.45609, 42.31711,
  62.93325, 61.13498, 56.34985, 54.50078, 54.76523, 55.36028, 56.07883,
    57.49861, 60.91235, 64.27374, 62.94181, 57.57324, 61.52948, 61.13857,
    59.22675, 57.33706, 58.14117, 59.95877, 62.03127, 61.85903, 63.29839,
    64.63973, 60.32702, 55.4477, 50.63879, 46.4235, 43.95219, 42.95353,
    42.48275, 42.33822,
  62.57624, 58.55171, 55.92805, 54.74291, 55.01993, 53.83324, 54.83759,
    55.92119, 60.71867, 62.87808, 56.08128, 52.13081, 55.11826, 56.10882,
    56.00755, 56.64916, 56.77021, 57.39772, 59.4935, 60.17274, 59.66681,
    60.30055, 62.23979, 61.63868, 55.43055, 47.8034, 44.32029, 43.55558,
    42.70387, 42.34908,
  63.40736, 62.24944, 58.62712, 58.01092, 61.01309, 62.45834, 61.45942,
    59.18478, 60.86362, 59.66646, 52.85073, 53.61496, 55.51146, 56.98595,
    56.63832, 58.04254, 58.50955, 56.11685, 55.78857, 55.78841, 54.91398,
    54.55742, 54.76465, 57.41684, 59.31456, 53.26657, 46.8224, 45.60381,
    44.25643, 42.52312,
  69.36842, 68.30103, 65.72414, 65.02837, 64.8601, 64.84222, 65.54134,
    66.59442, 68.27551, 65.71252, 57.31739, 59.60609, 61.58317, 63.5969,
    63.51203, 63.65428, 63.85379, 61.67469, 58.22012, 56.70961, 55.04271,
    53.94493, 53.64536, 53.88807, 56.78745, 59.49967, 54.89029, 48.06071,
    46.01223, 43.4967,
  70.68435, 68.91895, 62.97177, 61.31784, 63.04848, 63.45405, 64.14597,
    67.25246, 70.01759, 69.44304, 60.25675, 61.91073, 63.19474, 64.65945,
    65.00082, 66.6677, 66.69305, 66.30193, 63.6076, 60.0061, 57.87112,
    56.50154, 55.05138, 53.57558, 54.77345, 59.15765, 60.10612, 53.86214,
    49.67924, 45.9819,
  72.01112, 70.1912, 67.40459, 65.03239, 64.14175, 64.00175, 66.55254,
    69.16947, 70.26252, 67.76262, 66.04556, 65.89812, 66.22119, 65.29235,
    64.74008, 66.42091, 68.38739, 69.22116, 68.6524, 66.12668, 64.1998,
    62.9606, 59.85564, 57.01485, 57.29123, 58.50533, 60.93194, 56.18497,
    48.0673, 45.07823,
  71.6825, 69.91818, 67.34845, 65.19884, 64.76086, 62.79834, 66.56361,
    68.33377, 66.11755, 64.28782, 66.23805, 66.06443, 65.93724, 66.22392,
    67.21592, 68.62096, 70.47992, 70.81843, 70.53238, 70.08175, 69.42557,
    69.3829, 68.68323, 67.34697, 66.71506, 66.29008, 66.41151, 64.90058,
    51.19589, 43.02962,
  70.41541, 68.19437, 67.27893, 66.45126, 67.48738, 67.59814, 67.67433,
    66.60108, 60.88816, 62.68922, 63.84332, 64.29228, 65.06741, 66.15206,
    67.9907, 69.05819, 69.3021, 69.81325, 70.07638, 70.1226, 69.17531,
    67.8263, 65.02808, 64.59584, 65.48265, 65.90098, 65.75164, 65.94556,
    64.24413, 47.43212,
  63.97683, 63.83628, 64.28584, 64.74944, 66.47286, 68.11116, 67.46503,
    64.20444, 60.27121, 61.5424, 61.61346, 63.11357, 64.37672, 64.90293,
    65.58595, 65.69063, 64.61164, 63.31404, 59.95566, 56.14654, 54.89257,
    53.51037, 51.12798, 49.92841, 51.68376, 53.80492, 54.53622, 53.20414,
    53.15048, 48.71709,
  63.25124, 63.54769, 63.73789, 62.94332, 64.55247, 67.00751, 67.77849,
    65.32069, 60.66426, 64.25593, 65.409, 66.20792, 66.14692, 65.0461,
    64.18724, 63.00979, 57.39757, 51.92154, 50.87222, 49.29343, 47.23525,
    47.2961, 47.19961, 47.15686, 47.8677, 49.44939, 49.97834, 47.65964,
    44.67539, 42.34042,
  40.63199, 40.95095, 41.26019, 41.62635, 41.87302, 42.18886, 42.57191,
    43.02924, 43.53587, 44.15818, 45.66813, 45.70559, 43.69616, 44.13197,
    44.29868, 43.70254, 43.70215, 44.1295, 44.71188, 45.99683, 46.7317,
    46.17432, 46.81799, 48.12239, 48.73906, 48.26172, 51.17576, 51.32446,
    42.4257, 39.64445,
  46.4991, 47.14679, 47.10563, 48.08072, 48.24284, 48.5251, 49.2415,
    49.92683, 50.69498, 51.50046, 52.43593, 53.64071, 54.32044, 52.93583,
    52.01318, 52.04967, 50.88751, 51.04339, 51.89132, 52.60009, 52.36674,
    51.88721, 52.17159, 54.50757, 58.10862, 56.43669, 52.8521, 53.62474,
    43.68452, 40.73917,
  49.65808, 50.60321, 51.45074, 52.44705, 53.41684, 54.37735, 55.27041,
    56.34809, 57.50277, 58.51098, 59.45055, 60.63297, 61.73066, 63.12,
    63.54802, 61.88017, 61.44638, 61.644, 61.52385, 62.13803, 63.67264,
    65.04238, 64.94096, 65.0212, 66.2411, 64.02202, 58.75714, 52.93576,
    44.12292, 41.84996,
  55.40856, 57.09891, 58.82757, 60.66063, 62.40704, 63.6843, 63.96337,
    64.04803, 64.19032, 64.25144, 64.26215, 64.69025, 64.96613, 64.85979,
    65.73272, 66.72956, 66.97521, 66.69216, 66.84855, 67.48091, 68.3574,
    68.31745, 65.38604, 69.0037, 69.3089, 65.64417, 61.48845, 51.64644,
    44.0611, 40.39694,
  60.5878, 61.68515, 63.47185, 63.93655, 63.94373, 64.22375, 64.72939,
    64.95686, 65.111, 65.01722, 64.98856, 65.44447, 65.7737, 65.95264,
    66.27671, 67.06996, 67.49622, 66.80746, 66.09383, 68.47189, 68.73424,
    64.31555, 63.88622, 66.30669, 69.0998, 66.88295, 60.333, 59.88372,
    55.51181, 43.66707,
  64.0761, 64.46223, 64.89917, 65.10355, 64.70405, 64.76785, 65.48132,
    65.60833, 65.31843, 65.21443, 65.35363, 66.01661, 66.62538, 66.39317,
    66.61656, 67.95555, 69.53633, 69.21998, 68.19362, 68.31712, 66.36049,
    62.04865, 62.85139, 64.16363, 66.52943, 64.7794, 62.23076, 66.38413,
    64.0601, 42.39035,
  64.85859, 65.21638, 65.49945, 65.54671, 65.07935, 65.13495, 65.69701,
    65.7276, 65.26604, 65.12565, 65.1601, 65.14806, 65.05128, 65.19926,
    65.57661, 66.86784, 68.40488, 68.35438, 65.70605, 64.86832, 62.45932,
    60.95417, 61.63152, 63.99077, 63.71279, 60.0839, 62.54873, 66.5074,
    58.51594, 39.74657,
  65.02532, 65.28243, 65.47312, 65.53989, 65.0553, 64.96447, 65.38077,
    64.99152, 64.46597, 64.50768, 64.5852, 64.64533, 64.7001, 64.95435,
    65.50858, 66.70309, 68.17991, 68.187, 63.47956, 62.42954, 61.22066,
    61.20775, 63.21853, 64.50704, 61.36663, 59.88503, 66.03439, 64.23428,
    49.66211, 40.08457,
  66.72045, 67.00018, 67.22533, 67.08886, 66.57511, 66.68468, 66.85918,
    67.3434, 67.97681, 68.21437, 68.35935, 68.48451, 68.73578, 70.10968,
    71.00645, 70.06024, 71.04405, 72.21264, 72.17475, 70.9754, 70.11544,
    70.60338, 71.40928, 70.46085, 67.02762, 66.75156, 65.90684, 56.84232,
    43.4103, 39.72527,
  72.82047, 73.51331, 73.6143, 74.04206, 72.97496, 71.3215, 70.78923,
    71.59855, 72.03165, 72.68836, 73.1912, 73.91122, 73.68772, 72.57819,
    71.75672, 72.83995, 73.48037, 73.31772, 72.2486, 71.62666, 71.56143,
    70.67597, 69.39051, 63.84348, 66.92899, 68.71878, 62.76059, 44.53507,
    39.81907, 38.30282,
  74.19005, 74.62328, 76.22102, 76.19312, 77.42134, 76.33831, 75.15185,
    74.56307, 74.1757, 74.56075, 74.23714, 69.42127, 68.75932, 68.5283,
    68.92435, 69.72383, 70.54362, 70.50143, 69.46309, 66.44901, 67.35902,
    62.86793, 54.7572, 50.67762, 51.75112, 50.8115, 44.22416, 39.57468,
    39.11423, 38.25816,
  75.58242, 72.03923, 74.74333, 76.2258, 75.87843, 74.70263, 73.82754,
    71.07832, 68.1804, 67.86857, 67.13662, 65.92658, 66.12322, 66.66171,
    66.63554, 67.06167, 66.59163, 63.3932, 60.52599, 59.52739, 60.62058,
    56.27622, 48.9063, 53.77082, 55.91117, 44.54267, 39.48846, 40.11041,
    39.58811, 38.69835,
  80.99114, 81.03168, 82.29636, 82.98653, 81.96669, 78.72889, 71.70688,
    68.28098, 69.05329, 66.79062, 67.30157, 66.69637, 66.88783, 67.19473,
    66.72609, 66.7225, 67.67296, 64.63354, 61.85699, 62.79923, 60.8569,
    53.4653, 49.47835, 50.19405, 50.4638, 42.98153, 40.27187, 40.44786,
    40.44791, 39.24892,
  75.44588, 75.64488, 75.57175, 73.89521, 72.58911, 71.88789, 71.89574,
    72.42216, 70.05474, 69.8838, 70.59829, 68.96138, 70.01427, 70.51835,
    68.86473, 67.97253, 68.25538, 69.03902, 69.33469, 68.88166, 59.6961,
    53.24131, 52.58157, 45.53342, 42.18313, 41.34558, 40.01258, 39.44335,
    39.60181, 39.0438,
  68.53448, 68.42519, 68.20619, 67.8672, 67.89587, 69.17661, 72.96761,
    74.15821, 71.5816, 71.39645, 70.82867, 70.2584, 70.03878, 69.43279,
    68.67767, 67.75669, 68.12296, 68.88603, 69.83671, 68.25954, 54.69518,
    51.03794, 44.87347, 42.55942, 41.42765, 40.93268, 39.92496, 39.23291,
    38.8852, 38.55246,
  69.57951, 70.07951, 70.53376, 70.52734, 70.52223, 71.52789, 72.60218,
    72.4757, 71.90615, 71.08678, 70.48628, 68.96062, 68.06214, 68.41764,
    67.45649, 67.36277, 68.13863, 65.64991, 61.88025, 57.42259, 46.90355,
    45.86068, 43.29002, 42.31627, 41.64886, 40.82476, 39.89124, 39.33781,
    38.93721, 38.52136,
  69.45512, 69.45052, 69.59936, 69.78146, 70.42091, 70.49265, 71.05286,
    71.74415, 71.31966, 70.60299, 69.29748, 69.41625, 70.21886, 68.46624,
    67.23502, 67.19743, 67.20802, 61.14677, 61.01064, 58.2485, 45.64573,
    45.76133, 43.73881, 42.37793, 41.32346, 40.8668, 39.78841, 38.87004,
    38.69653, 38.48089,
  67.80491, 68.28882, 68.27492, 68.64737, 68.8247, 69.30174, 69.55524,
    69.98405, 70.44145, 69.5779, 69.624, 69.9778, 69.08403, 68.25774,
    68.0415, 67.26597, 62.21513, 56.99998, 58.98338, 55.33919, 45.90348,
    44.9693, 43.19649, 41.98473, 40.36814, 39.94156, 39.50156, 38.58676,
    38.45054, 38.3134,
  69.89771, 68.88418, 67.60612, 66.94447, 67.45203, 67.50752, 67.95667,
    68.52272, 68.36106, 68.29138, 68.7798, 68.17493, 66.90335, 67.39999,
    67.85606, 69.01692, 71.07039, 72.50087, 72.60625, 66.45966, 53.91002,
    46.48691, 42.99162, 41.78845, 39.93243, 39.37299, 39.10207, 38.59962,
    38.40847, 38.29328,
  69.56461, 68.3609, 67.1589, 66.45654, 66.99406, 67.37919, 67.78643,
    68.09756, 68.35308, 69.02039, 69.02349, 67.64678, 67.55672, 67.69788,
    68.09071, 69.06091, 70.58106, 69.66148, 68.11423, 65.41293, 58.13932,
    49.86612, 44.05471, 42.44759, 40.72516, 39.5785, 39.09748, 38.66617,
    38.40075, 38.30495,
  68.9203, 67.994, 66.69324, 66.08298, 66.47722, 66.76101, 67.11704,
    67.41128, 67.71986, 68.1049, 67.4142, 66.33392, 66.50088, 66.54283,
    66.55949, 62.62678, 60.1455, 58.64436, 58.49418, 57.23111, 55.16307,
    52.96848, 48.35263, 44.5043, 41.82072, 40.18459, 39.08876, 38.66862,
    38.42627, 38.3227,
  69.10341, 67.48559, 66.27406, 65.48075, 65.72157, 65.68454, 65.87106,
    65.97578, 66.45145, 66.43239, 64.80807, 62.13168, 62.51235, 61.19092,
    58.95206, 56.68663, 54.33789, 52.76482, 52.12436, 51.263, 51.82416,
    52.4232, 51.06158, 49.87499, 45.42249, 41.20415, 39.26784, 38.93122,
    38.48788, 38.31466,
  68.7639, 67.39565, 65.87106, 64.97699, 65.36012, 65.42754, 65.09524,
    64.65068, 64.84225, 62.72101, 58.39919, 58.45688, 58.70126, 58.12312,
    56.41368, 55.14756, 53.39452, 50.59092, 49.19121, 48.54581, 49.18564,
    49.82506, 48.04802, 48.34504, 47.90132, 43.56293, 40.11728, 39.83584,
    39.07061, 38.39003,
  70.33287, 69.09955, 68.03255, 67.33072, 67.32217, 67.08524, 67.17419,
    67.43295, 67.86371, 65.39994, 61.22433, 62.81638, 63.23448, 62.7501,
    60.83329, 58.42216, 56.23486, 53.26802, 50.12077, 49.10925, 49.32887,
    48.90926, 47.36174, 46.37009, 46.53955, 46.36345, 43.17841, 40.57602,
    39.76252, 38.73282,
  72.11685, 72.54937, 70.0844, 69.08539, 69.25397, 69.14269, 69.09763,
    69.61372, 70.59207, 69.75327, 64.98651, 66.41388, 66.41486, 64.99342,
    62.42761, 59.88512, 56.79325, 54.39753, 51.43766, 48.95354, 48.76209,
    48.31128, 46.8405, 45.57328, 44.63268, 45.59095, 45.63503, 42.96856,
    41.39683, 39.78656,
  74.71165, 75.4698, 73.52733, 72.03308, 71.48147, 71.0749, 71.59688,
    72.33598, 72.11318, 69.84215, 68.02824, 68.42101, 67.92244, 64.79079,
    60.95727, 58.40397, 56.03012, 54.0815, 51.94443, 49.69488, 49.53589,
    49.2489, 47.06668, 45.27127, 44.82963, 45.04573, 46.02276, 44.35775,
    41.03843, 39.52025,
  75.33853, 75.76952, 73.68055, 72.41273, 72.29995, 71.78413, 72.12543,
    72.34955, 71.0737, 68.39124, 68.35634, 68.30621, 67.17682, 64.42088,
    61.60449, 58.9662, 56.80405, 55.67998, 54.33609, 53.1054, 54.37867,
    56.15984, 54.99691, 51.44513, 49.16906, 48.4445, 49.18392, 47.83496,
    41.69609, 38.52403,
  75.34422, 75.45676, 74.04237, 73.54177, 74.06163, 73.77751, 73.23196,
    72.4974, 70.41654, 70.33177, 70.27731, 70.49324, 69.85793, 68.00992,
    66.4223, 64.02949, 61.4312, 60.39175, 59.88207, 59.62751, 59.93007,
    58.44919, 54.77549, 52.15435, 50.51558, 49.77655, 48.91297, 50.21176,
    47.39818, 40.32489,
  71.33922, 71.50886, 72.56497, 73.3535, 73.88609, 74.31208, 73.32822,
    71.35676, 70.5106, 70.39159, 69.96208, 69.58284, 69.35532, 69.56385,
    70.26861, 68.57958, 65.72059, 63.26286, 59.57116, 55.76619, 54.07212,
    52.01617, 49.54778, 47.79456, 47.30539, 47.03917, 46.13821, 44.54366,
    44.03707, 41.32807,
  69.76984, 70.00195, 70.50515, 70.67561, 71.41143, 72.55622, 72.42315,
    70.43189, 69.18315, 69.30031, 69.28683, 69.04163, 68.58848, 68.21955,
    68.28008, 64.5556, 58.66743, 53.49213, 51.03573, 48.65538, 46.71141,
    45.82248, 44.99413, 44.21066, 43.72557, 43.7076, 43.16944, 41.59478,
    39.92519, 38.52939,
  34.80149, 34.89823, 34.97809, 35.05098, 35.07703, 35.141, 35.2284,
    35.37298, 35.56712, 35.80266, 36.76288, 36.91265, 35.52273, 35.71806,
    35.87078, 35.47781, 35.45231, 35.68241, 35.93932, 36.74847, 37.285,
    36.79733, 36.99925, 37.94226, 38.66214, 38.50664, 41.1513, 42.53417,
    37.23783, 35.48423,
  36.49709, 36.69647, 36.45083, 36.85736, 36.72064, 36.64385, 36.83956,
    37.05562, 37.29486, 37.55996, 37.95804, 38.59343, 39.04668, 38.11473,
    37.50312, 37.73826, 37.26047, 37.64036, 38.45782, 39.26508, 39.49627,
    39.4435, 39.99815, 41.47962, 46.14732, 47.15427, 41.87116, 44.09338,
    37.98897, 36.13381,
  37.95358, 38.15156, 38.25631, 38.45029, 38.59553, 38.76171, 38.94591,
    39.18675, 39.45493, 39.69525, 40.00699, 40.58081, 40.98872, 41.5644,
    41.78247, 40.8243, 40.98621, 41.81587, 42.37224, 43.31961, 45.02314,
    47.04797, 48.06173, 47.47038, 51.40095, 53.55874, 45.11322, 43.33215,
    38.01039, 36.81765,
  41.2968, 41.76944, 42.33765, 42.96677, 43.60552, 44.43331, 44.69489,
    44.60141, 44.90576, 45.44652, 45.68829, 46.16433, 46.15888, 45.5125,
    46.57787, 47.57094, 46.5887, 45.39804, 46.27361, 47.40613, 50.015,
    50.91835, 48.85637, 53.52767, 55.64023, 48.93898, 47.78106, 42.32161,
    38.00056, 35.92557,
  46.33225, 46.52198, 47.21844, 47.93988, 48.3959, 48.67071, 48.8456,
    48.97852, 49.71032, 50.32416, 50.15284, 50.35062, 50.39801, 50.4475,
    50.38918, 50.36938, 49.23767, 47.60522, 47.79038, 52.77428, 54.6922,
    46.75397, 46.76735, 48.23729, 49.9626, 48.73989, 44.92174, 44.92308,
    44.30152, 38.14487,
  50.26377, 51.11847, 52.2359, 53.63408, 53.57589, 53.20338, 53.89465,
    54.29645, 54.36847, 55.09776, 56.05843, 58.47914, 60.88812, 59.8382,
    58.33474, 66.14521, 73.98344, 60.41784, 50.44196, 51.06169, 48.47402,
    45.01655, 45.82864, 47.04036, 49.36067, 47.98969, 50.96491, 66.5808,
    58.07034, 36.93068,
  55.25586, 56.79143, 58.2918, 60.06387, 60.7849, 61.37037, 63.00087,
    64.87035, 64.65166, 63.75254, 63.27187, 61.22858, 58.14408, 57.15784,
    60.90931, 66.18306, 60.35096, 52.01625, 48.29101, 47.68382, 46.12761,
    45.2543, 45.95519, 48.35139, 49.12114, 45.37365, 54.89248, 71.68658,
    55.15458, 35.12048,
  60.83222, 62.60331, 64.16215, 65.58583, 65.18896, 66.38808, 67.36588,
    62.75515, 58.96906, 57.79784, 56.12399, 54.13855, 52.26365, 51.50963,
    51.35748, 51.17625, 50.32201, 49.01692, 46.2541, 45.64286, 44.83182,
    44.69744, 46.26772, 48.16682, 46.97196, 44.63562, 55.50164, 60.64124,
    42.02661, 35.80409,
  65.11925, 65.46942, 65.87184, 65.15874, 63.47414, 63.01237, 59.68485,
    57.17811, 56.87707, 56.35099, 55.45042, 54.50761, 53.91188, 56.924,
    58.39972, 52.30383, 51.01609, 52.21622, 51.65501, 48.47427, 46.20857,
    48.49413, 52.88356, 52.83165, 47.86303, 48.18147, 51.20447, 47.69949,
    38.06186, 35.65386,
  69.03096, 69.44178, 69.69994, 69.89579, 69.33633, 63.54489, 57.87745,
    59.12401, 59.5913, 61.24763, 63.25835, 66.44603, 66.09355, 62.24842,
    57.79193, 57.91627, 58.12905, 57.3555, 55.07903, 53.57924, 53.99527,
    53.46339, 52.56347, 48.64933, 56.06311, 69.28603, 55.13195, 38.9196,
    35.91991, 34.65092,
  72.44817, 72.22469, 72.6085, 71.93968, 71.74673, 71.5262, 70.95585,
    71.09087, 71.44672, 73.16193, 74.49679, 64.98659, 59.78378, 58.26469,
    57.10574, 56.6641, 56.65049, 55.62516, 53.88506, 52.83448, 54.48975,
    52.23206, 46.73058, 43.16611, 45.00901, 46.3499, 40.25882, 35.59289,
    35.14251, 34.546,
  78.04979, 74.16331, 77.58286, 78.66377, 78.30782, 76.92078, 75.79482,
    72.65565, 69.60593, 69.95741, 69.4635, 61.61155, 62.93136, 62.03061,
    56.3805, 55.30877, 52.88461, 51.47106, 49.78256, 49.05345, 50.27741,
    47.76934, 41.62597, 45.83351, 48.30154, 38.28156, 35.27568, 35.67417,
    35.42532, 34.82932,
  84.92533, 85.15051, 87.659, 87.91318, 86.49548, 82.25513, 74.30482,
    69.87073, 70.12947, 68.49662, 68.73187, 68.4952, 69.17242, 69.26225,
    59.14727, 53.5811, 51.39273, 49.62416, 47.95094, 49.02565, 48.88708,
    44.44574, 40.85125, 44.31233, 46.07262, 37.24823, 35.75502, 35.90983,
    35.99493, 35.21249,
  82.01323, 83.93903, 82.94404, 80.33537, 77.66421, 75.80231, 75.01635,
    74.76541, 72.27142, 71.28854, 72.21669, 71.00634, 72.19217, 73.02723,
    72.61417, 63.31508, 52.21447, 53.23215, 53.32553, 52.13501, 46.98578,
    45.74243, 48.47916, 40.89279, 37.67543, 36.63038, 35.77852, 35.3715,
    35.53591, 35.11603,
  73.54202, 73.03147, 72.05398, 70.81571, 69.83437, 71.56353, 77.01177,
    76.97192, 73.4937, 72.8168, 71.61137, 70.12801, 69.81413, 71.17429,
    72.36157, 58.31727, 56.32066, 53.8804, 54.4035, 55.39307, 51.3758,
    44.84243, 39.35929, 37.33184, 36.52297, 36.52246, 35.7776, 35.23281,
    35.02356, 34.78171,
  70.03408, 70.08576, 70.30316, 70.07498, 69.93045, 70.69885, 71.56183,
    71.20456, 70.34985, 69.46463, 69.10885, 68.12129, 63.77598, 63.68428,
    59.30748, 55.26458, 53.56249, 49.74461, 48.49554, 46.98674, 40.89034,
    39.10743, 37.10439, 36.67915, 36.67076, 36.35921, 35.77705, 35.31225,
    35.00913, 34.73033,
  69.265, 69.33747, 69.42757, 69.41169, 69.63676, 69.17521, 69.22517,
    69.75667, 69.38251, 68.77934, 65.22444, 64.64548, 66.41833, 60.61608,
    55.51167, 52.09346, 49.0399, 46.03492, 46.82705, 45.75355, 38.2538,
    38.53887, 37.58665, 36.74951, 36.38356, 36.34869, 35.70226, 35.04238,
    34.88022, 34.7109,
  68.31744, 68.75588, 68.5907, 68.61751, 68.32722, 67.82179, 67.22448,
    66.7631, 66.41756, 63.639, 63.71832, 64.95648, 61.80235, 58.8024,
    57.32079, 51.63094, 45.71633, 42.81659, 45.14021, 44.0496, 38.43412,
    38.36424, 37.58129, 36.88431, 35.96827, 35.82145, 35.50185, 34.84806,
    34.72321, 34.61537,
  69.7477, 68.63989, 65.31112, 63.15515, 62.39952, 61.39735, 60.96621,
    60.85148, 59.71258, 58.66489, 59.73117, 57.67081, 52.04607, 51.3918,
    50.46732, 48.64538, 48.66834, 49.33056, 51.53992, 50.48288, 44.27582,
    39.83118, 37.47492, 36.92899, 35.76637, 35.41481, 35.23606, 34.83932,
    34.69017, 34.59657,
  66.20227, 64.15396, 61.10636, 58.51639, 57.72342, 57.01978, 56.44775,
    55.87994, 55.38519, 56.82882, 56.62941, 51.88148, 50.1212, 49.54077,
    48.64782, 47.66734, 48.51898, 49.88177, 50.63266, 50.46836, 46.88705,
    41.69682, 37.81931, 37.19566, 36.21766, 35.48735, 35.18216, 34.87801,
    34.6929, 34.60508,
  62.31487, 60.52534, 57.6288, 55.35288, 54.44687, 53.90399, 53.45698,
    53.17721, 53.615, 55.12397, 53.46164, 50.13343, 50.63826, 50.05445,
    48.41759, 46.46789, 45.64988, 45.09392, 45.09442, 44.4116, 43.0914,
    42.0727, 40.07167, 38.22389, 36.80534, 35.84701, 35.19621, 34.88064,
    34.69971, 34.62377,
  61.56601, 58.62172, 56.21461, 54.55207, 53.75111, 52.78866, 52.68123,
    52.47768, 53.87554, 54.47178, 51.37659, 49.19697, 49.0118, 47.49827,
    45.46705, 43.8546, 42.47297, 41.50999, 41.07932, 40.34513, 41.56824,
    42.58165, 40.82276, 41.15302, 38.86724, 36.44446, 35.27643, 35.02742,
    34.74021, 34.61843,
  60.42304, 58.63248, 56.0538, 54.61559, 54.95129, 54.9433, 54.04939,
    52.58722, 52.74525, 51.4927, 48.03238, 47.0346, 46.18305, 44.78074,
    42.92859, 42.16429, 41.59483, 40.21038, 39.52314, 39.05798, 40.24778,
    41.05698, 38.83414, 39.9128, 40.12151, 37.68958, 35.6829, 35.57263,
    35.10892, 34.66422,
  60.77006, 59.45836, 58.20118, 57.43247, 56.81865, 55.74949, 55.29924,
    54.44395, 54.16991, 50.6667, 46.74584, 46.69355, 46.17591, 45.29282,
    43.944, 42.955, 42.5458, 41.46595, 39.80326, 39.1008, 39.1721, 39.07694,
    38.37097, 38.23434, 38.91035, 39.21359, 37.50663, 35.98427, 35.52362,
    34.87433,
  60.39951, 60.53268, 57.51294, 56.10476, 55.84254, 54.93488, 53.52932,
    52.82159, 53.61675, 50.89342, 46.73359, 47.05942, 46.83698, 45.85601,
    44.54306, 43.76947, 42.78529, 42.10513, 40.80091, 39.341, 39.21951,
    39.22884, 38.80777, 38.05293, 37.51405, 38.61517, 38.84156, 37.27013,
    36.5012, 35.50121,
  61.20102, 62.44807, 60.58646, 57.81839, 55.78827, 54.38989, 54.70738,
    55.11148, 53.11871, 49.99292, 48.19187, 48.29462, 48.06624, 46.21252,
    44.06774, 43.15959, 42.49991, 42.01224, 41.14384, 39.74833, 39.66842,
    39.7327, 38.59449, 37.67377, 37.63604, 38.07321, 39.09973, 38.26832,
    36.36331, 35.33669,
  62.09654, 62.38372, 59.00016, 56.69993, 55.51047, 54.07135, 54.72642,
    54.3129, 51.21177, 48.98321, 48.73219, 48.53863, 47.61141, 45.61808,
    43.86567, 42.685, 41.89235, 41.6599, 41.04771, 39.96806, 40.49665,
    42.0112, 42.15187, 40.73474, 39.91711, 39.84198, 40.92738, 40.46482,
    36.69117, 34.71875,
  61.46976, 60.4663, 58.10624, 57.22957, 56.91028, 55.64725, 54.96354,
    52.79747, 49.18773, 48.52954, 48.08989, 47.7226, 46.78559, 45.21756,
    44.27368, 43.35808, 42.46581, 42.4754, 42.8321, 43.06145, 43.78244,
    43.84687, 42.49986, 41.31463, 40.68664, 40.60318, 40.44086, 41.76429,
    40.19732, 35.82691,
  59.07259, 57.61877, 57.76019, 58.20393, 57.94831, 57.96623, 55.55839,
    50.71746, 48.14814, 47.94505, 46.9619, 46.27162, 45.75168, 45.52269,
    45.81618, 45.89208, 45.79047, 45.90484, 44.77238, 43.0161, 42.49066,
    41.63983, 40.35187, 39.50495, 39.41858, 39.55666, 39.28039, 38.56473,
    38.54251, 36.57112,
  58.1465, 57.74971, 57.18324, 56.11179, 55.77768, 57.47116, 57.40847,
    52.31028, 49.1689, 49.9817, 50.50803, 50.78102, 50.31596, 49.55871,
    48.69592, 47.59362, 45.60896, 43.35009, 42.09067, 40.67079, 39.56665,
    39.03503, 38.5529, 38.14957, 37.92428, 38.03788, 37.74468, 36.81443,
    35.87716, 34.86335,
  31.70529, 31.76044, 31.80197, 31.82689, 31.82747, 31.83877, 31.86264,
    31.92914, 32.05572, 32.19078, 32.96728, 33.12942, 32.06264, 32.20893,
    32.34638, 32.01454, 31.92947, 32.02315, 32.11588, 32.66648, 32.99334,
    32.4922, 32.48026, 33.11608, 33.59217, 33.40894, 35.66257, 37.1756,
    33.59683, 32.34336,
  32.30276, 32.41968, 32.18022, 32.45169, 32.31912, 32.19443, 32.29966,
    32.41257, 32.55778, 32.74921, 33.07624, 33.59237, 33.93602, 33.25575,
    32.80636, 32.94251, 32.48818, 32.6367, 33.16813, 33.69497, 33.72362,
    33.4465, 33.76339, 34.73067, 38.92108, 40.46112, 36.20112, 38.54877,
    34.21223, 32.80938,
  32.41045, 32.44066, 32.43673, 32.50283, 32.51406, 32.54218, 32.60999,
    32.71954, 32.844, 32.97095, 33.11179, 33.51506, 33.82546, 34.29435,
    34.52816, 33.81207, 33.85056, 34.39675, 34.68111, 35.22452, 36.40198,
    37.94059, 39.05045, 38.67105, 43.22948, 46.44773, 38.51279, 38.08229,
    34.17876, 33.3428,
  33.02125, 33.12157, 33.40786, 33.69666, 34.01102, 34.54949, 34.69143,
    34.49669, 34.63848, 34.96194, 35.08572, 35.403, 35.41125, 35.09076,
    36.18737, 37.32749, 36.88742, 36.08411, 36.78953, 37.68727, 40.0153,
    41.31024, 39.89033, 44.68331, 47.3825, 41.36217, 40.89154, 37.28713,
    34.14314, 32.70714,
  34.77677, 34.69852, 35.14917, 35.62218, 35.95941, 36.13648, 36.23035,
    36.25254, 36.76641, 37.16196, 36.91136, 36.98502, 37.10584, 37.52739,
    38.24917, 38.96732, 38.52035, 38.00996, 38.54553, 43.26149, 45.47026,
    38.96972, 38.89009, 40.35194, 41.94413, 40.86367, 38.29359, 38.11929,
    38.32871, 34.35809,
  36.45748, 36.93835, 37.75607, 38.7792, 38.6492, 38.19206, 38.57038,
    38.75457, 38.70094, 39.15905, 39.72368, 41.65229, 43.90442, 43.92398,
    43.09002, 51.67154, 61.93534, 49.51132, 41.47872, 42.65593, 40.83438,
    37.63425, 38.06768, 38.78831, 40.7735, 39.87673, 42.84639, 57.15893,
    51.13389, 33.52996,
  38.64395, 39.47568, 40.50756, 41.70354, 42.12561, 42.50692, 43.97145,
    45.96085, 46.55639, 46.64987, 47.08431, 46.30786, 44.575, 44.12512,
    49.29476, 57.39376, 52.66937, 43.46444, 40.45472, 39.88652, 38.4721,
    37.66114, 38.14437, 40.01786, 41.11795, 38.05186, 47.83173, 65.56301,
    50.52859, 32.04984,
  41.7709, 43.13581, 44.70153, 46.37507, 46.84072, 48.77038, 50.90433,
    48.72058, 46.70609, 46.41264, 45.48891, 43.91946, 42.2836, 41.71376,
    42.48619, 43.31361, 42.14461, 40.82087, 38.81851, 38.35201, 37.68689,
    37.4608, 38.65379, 40.28138, 39.79501, 37.5126, 49.84217, 56.90966,
    37.93446, 33.00643,
  47.35842, 48.48286, 49.71294, 50.16315, 49.91255, 50.62061, 48.74701,
    46.88057, 46.53819, 45.90359, 44.7305, 43.31799, 42.32559, 44.67515,
    46.16122, 41.9212, 41.34781, 42.57329, 42.28823, 39.92329, 37.9867,
    39.52162, 43.08238, 43.32783, 39.60285, 39.95987, 44.23806, 43.03974,
    35.23079, 32.93718,
  53.27629, 55.47329, 55.90036, 56.35241, 54.73933, 50.4413, 45.6404,
    45.7671, 45.46242, 45.7514, 46.83836, 49.75522, 49.93147, 47.60016,
    44.64278, 44.63377, 45.11138, 44.8669, 43.5584, 43.0541, 43.50599,
    43.83688, 44.02885, 41.52019, 48.20272, 59.787, 49.06211, 35.76648,
    33.30775, 31.87716,
  74.80477, 74.26254, 71.00948, 61.15672, 58.94344, 55.79982, 51.90158,
    53.87619, 55.26582, 63.98586, 71.41831, 50.18038, 44.74185, 43.55414,
    42.67289, 43.15777, 44.65688, 44.30975, 43.14425, 42.79519, 45.35176,
    44.53536, 40.48845, 37.69154, 40.79567, 43.68506, 37.82326, 32.81738,
    32.30728, 31.73495,
  78.48547, 73.69265, 76.40384, 77.75505, 78.34227, 71.95376, 71.34695,
    64.51881, 54.07065, 57.1539, 56.30516, 44.297, 45.8657, 46.1763,
    42.39153, 43.37766, 42.29678, 41.84737, 40.93416, 41.01946, 43.58971,
    42.02476, 36.72935, 40.38107, 42.60635, 34.94205, 32.26291, 32.66106,
    32.54604, 31.98089,
  81.53716, 81.6291, 86.21647, 87.88151, 88.65005, 85.93157, 78.57028,
    56.95841, 56.50526, 52.68077, 51.57283, 46.16893, 49.67008, 50.76459,
    44.13231, 43.15995, 42.44463, 41.3241, 40.07566, 41.93394, 43.14827,
    39.31675, 36.0599, 40.39942, 42.13712, 33.98659, 32.58952, 32.83149,
    33.04418, 32.30936,
  83.0548, 87.70317, 87.27136, 85.53059, 82.78111, 79.8615, 77.09404,
    76.17135, 75.39529, 72.24738, 76.55733, 76.35017, 76.13722, 73.89325,
    63.35863, 50.99466, 42.62745, 44.24175, 45.25858, 45.63935, 41.81856,
    40.6794, 43.08977, 37.48409, 34.70226, 33.35484, 32.63394, 32.34713,
    32.66229, 32.25182,
  78.16438, 78.3147, 74.88578, 70.67781, 66.29102, 74.40112, 79.46793,
    79.87936, 76.88631, 76.82001, 76.79724, 64.67747, 53.05103, 58.26436,
    62.62495, 46.87401, 46.58907, 45.93277, 48.79166, 50.32573, 45.21949,
    40.53808, 36.37199, 34.0389, 33.14064, 33.41467, 32.73832, 32.27416,
    32.15574, 31.92804,
  65.13531, 62.94071, 61.87491, 60.85028, 61.3939, 65.83355, 70.42087,
    67.59419, 64.16216, 60.74361, 56.15762, 49.90437, 46.97567, 49.35498,
    48.34562, 45.71347, 46.33564, 43.98848, 44.41125, 43.95506, 37.73946,
    35.30828, 33.37999, 33.19737, 33.48262, 33.32776, 32.80532, 32.3726,
    32.11837, 31.86283,
  60.61685, 58.88363, 58.04184, 57.80166, 58.13246, 57.57905, 56.61929,
    55.86975, 54.11539, 51.72146, 47.89521, 48.56795, 52.23325, 48.86765,
    45.73977, 44.7389, 43.23512, 40.89352, 42.7147, 42.02907, 34.27319,
    34.48907, 33.96894, 33.35315, 33.18781, 33.32368, 32.76393, 32.11761,
    31.99813, 31.85357,
  56.62901, 56.18788, 55.00483, 54.39622, 53.36686, 52.65504, 52.08138,
    51.5633, 50.60746, 48.58238, 48.66553, 51.12143, 49.69271, 48.27101,
    49.11572, 45.62638, 40.57108, 37.77507, 40.8902, 40.32783, 34.55848,
    34.74323, 34.27541, 33.675, 32.82651, 32.85216, 32.56287, 31.94014,
    31.84371, 31.76779,
  56.04359, 54.80888, 52.16348, 50.25599, 49.46264, 48.60913, 48.21933,
    48.17352, 47.28479, 46.51633, 48.25586, 47.19871, 42.11309, 42.09622,
    42.38784, 41.24686, 41.2263, 41.74852, 44.68906, 44.31332, 38.75013,
    35.84605, 34.44452, 33.85412, 32.7365, 32.46701, 32.31209, 31.93573,
    31.79839, 31.73775,
  53.68413, 52.02488, 49.52772, 47.45365, 46.89308, 46.40735, 46.02396,
    45.63239, 45.16095, 46.61633, 46.62276, 41.60936, 39.08851, 38.89537,
    38.65728, 38.0873, 39.52936, 41.57609, 43.57338, 44.65926, 41.86274,
    37.78212, 34.80283, 34.06576, 33.15421, 32.52228, 32.24446, 31.96443,
    31.8066, 31.73987,
  50.93952, 50.12172, 47.74979, 45.86536, 45.13015, 44.6586, 44.09435,
    43.46505, 43.47184, 44.75391, 42.48096, 38.19871, 38.48122, 38.79084,
    38.47853, 37.69525, 37.81147, 38.13984, 39.21543, 39.61227, 38.94741,
    38.34631, 36.79917, 34.93122, 33.5979, 32.82516, 32.25592, 31.97055,
    31.82481, 31.74863,
  49.65871, 48.32383, 46.23431, 44.80526, 43.95124, 42.75843, 42.25624,
    41.70221, 42.8804, 43.35713, 39.8896, 37.56309, 38.12659, 38.10504,
    37.67222, 37.21901, 36.55929, 36.11618, 36.11975, 35.70306, 36.98549,
    38.04593, 37.50396, 38.05833, 35.86739, 33.48318, 32.36017, 32.12583,
    31.86811, 31.76515,
  48.48268, 46.90828, 44.5429, 43.13609, 43.39081, 43.44852, 42.84287,
    41.85973, 42.74521, 41.89428, 38.32144, 37.45308, 37.44896, 37.26071,
    36.61018, 36.67635, 36.48452, 35.30632, 34.76395, 34.54175, 35.88273,
    36.54486, 35.23351, 36.8541, 37.21875, 34.6578, 32.67185, 32.62624,
    32.20246, 31.81399,
  47.421, 45.88611, 44.87005, 44.40419, 44.34002, 44.09191, 44.54184,
    44.74157, 45.52503, 42.39877, 38.08162, 37.85293, 37.80352, 37.89844,
    37.55959, 37.3011, 37.39763, 36.53222, 35.06778, 34.67109, 35.03502,
    35.03998, 34.54356, 34.75805, 35.85331, 36.21912, 34.43464, 33.01607,
    32.59204, 31.98849,
  46.8748, 47.32407, 44.83764, 44.00918, 44.45359, 44.38202, 43.8566,
    44.01699, 45.59646, 42.71832, 37.95602, 37.883, 38.07026, 38.06478,
    37.87031, 37.89666, 37.51438, 37.26059, 36.01045, 34.62548, 34.83599,
    35.12552, 34.94962, 34.27114, 33.80748, 35.1146, 35.41208, 33.99908,
    33.47738, 32.53152,
  47.93799, 49.62696, 48.3414, 46.34715, 44.88197, 43.83981, 44.74919,
    45.97408, 44.52842, 41.14932, 38.60685, 38.52682, 38.93581, 38.24862,
    37.30231, 37.25436, 37.10449, 37.08118, 36.35347, 34.93981, 35.29255,
    35.69167, 34.61519, 33.73014, 33.63553, 34.20643, 35.51187, 34.85465,
    33.35924, 32.39169,
  49.27615, 50.23632, 47.23069, 45.26924, 44.30215, 43.21042, 44.52004,
    45.07722, 42.14842, 39.54824, 38.87996, 38.81226, 38.66635, 37.81467,
    37.19905, 36.87051, 36.58438, 36.70288, 36.13612, 34.87391, 35.62472,
    37.43769, 37.70873, 36.25437, 35.42084, 35.55881, 37.12477, 37.01029,
    33.58378, 31.79101,
  48.63671, 48.13774, 46.01069, 45.28036, 45.40596, 44.75889, 45.04494,
    43.54415, 39.99263, 39.1466, 38.55241, 38.35379, 38.11299, 37.53411,
    37.58405, 37.27341, 36.54628, 36.61954, 36.83688, 36.81337, 38.19437,
    39.00901, 37.92405, 36.59451, 35.90505, 36.07533, 36.30194, 38.16978,
    36.78899, 32.76723,
  45.93164, 44.71284, 45.0657, 46.11757, 46.82242, 47.82251, 46.22669,
    42.02347, 39.49097, 39.06177, 37.65483, 36.64336, 36.28798, 36.71937,
    37.82317, 38.41037, 38.62102, 39.1675, 38.27941, 36.75857, 36.8212,
    36.4141, 35.30245, 34.59998, 34.72715, 35.1511, 35.2043, 35.00355,
    35.47592, 33.4851,
  45.00865, 44.95284, 44.80086, 44.33699, 44.57328, 47.06877, 47.70108,
    42.79418, 39.50595, 39.71907, 39.60184, 39.52883, 39.38737, 39.86754,
    40.46848, 40.37608, 39.19176, 37.5655, 36.56885, 35.31075, 34.54762,
    34.23547, 33.98612, 33.77198, 33.78487, 34.1912, 34.21775, 33.57758,
    32.90718, 32.03236,
  25.22817, 25.25784, 25.29526, 25.33168, 25.32068, 25.31923, 25.33152,
    25.37239, 25.44371, 25.54642, 26.42269, 26.58342, 25.52899, 25.69673,
    25.82521, 25.47393, 25.38373, 25.42883, 25.4647, 26.02719, 26.34512,
    25.81954, 25.76365, 26.32738, 26.64743, 26.31473, 28.80029, 30.6125,
    27.26118, 25.97797,
  25.67015, 25.75136, 25.49555, 25.77234, 25.62203, 25.4607, 25.53573,
    25.61278, 25.72943, 25.89606, 26.27761, 26.86522, 27.21577, 26.51863,
    26.10584, 26.17351, 25.65472, 25.72486, 26.20197, 26.71491, 26.68387,
    26.19892, 26.26201, 27.15898, 31.16899, 32.13605, 29.3085, 32.47263,
    28.05102, 26.5553,
  25.60645, 25.6362, 25.61672, 25.65534, 25.62543, 25.61369, 25.64245,
    25.73621, 25.83654, 25.90238, 26.02518, 26.44891, 26.7659, 27.23771,
    27.38416, 26.53355, 26.43445, 26.84802, 26.93632, 27.2459, 28.17801,
    29.62684, 30.65506, 30.30112, 34.93619, 37.82389, 31.72515, 31.9965,
    27.93544, 27.11259,
  25.78445, 25.82214, 26.02091, 26.21381, 26.50017, 27.01855, 27.08634,
    26.82251, 26.89097, 27.16832, 27.26649, 27.58966, 27.46243, 27.05823,
    28.10594, 29.15524, 28.51333, 27.46314, 27.80942, 28.40269, 30.96544,
    32.43483, 31.27611, 35.89838, 38.09571, 33.99454, 34.48193, 31.35017,
    27.93079, 26.39677,
  26.76349, 26.52295, 26.83608, 27.20733, 27.52424, 27.71569, 27.6915,
    27.56921, 28.09993, 28.48802, 28.19319, 28.1245, 28.02767, 28.35309,
    29.11237, 29.74499, 29.07018, 28.36294, 28.94159, 33.62031, 35.56548,
    30.27926, 30.13524, 32.0165, 33.88519, 33.26808, 31.43253, 31.68647,
    32.41964, 28.17556,
  27.62064, 27.83133, 28.56319, 29.58932, 29.49278, 28.93581, 29.0694,
    28.93761, 28.57301, 28.65557, 28.76564, 30.553, 32.87055, 32.95982,
    32.42588, 39.87394, 47.94262, 38.59981, 32.22085, 34.03392, 32.3191,
    28.84329, 29.29328, 30.17143, 32.68274, 32.22935, 34.53988, 47.72663,
    43.792, 27.55825,
  29.10696, 29.55822, 30.34476, 31.29517, 31.45048, 31.31928, 32.28502,
    34.00624, 34.3084, 34.14793, 34.61958, 34.10703, 32.81649, 32.93347,
    38.19516, 45.74779, 42.7477, 34.68187, 31.73387, 31.34309, 29.78545,
    28.76991, 29.27023, 31.6439, 33.20124, 30.56992, 39.89894, 56.38186,
    43.72951, 26.01313,
  30.99035, 31.66281, 32.77858, 34.025, 34.14146, 36.26151, 38.81205,
    36.77559, 34.90176, 34.74039, 34.10684, 32.68547, 31.31481, 31.28555,
    33.08644, 34.61589, 33.46128, 32.03598, 30.08035, 29.64221, 28.96759,
    28.68249, 30.02458, 32.37487, 32.10046, 30.29185, 42.72102, 49.27157,
    32.48968, 26.34008,
  34.76271, 35.45395, 36.75809, 37.3279, 37.6828, 39.39981, 38.3126,
    36.57806, 36.27687, 35.66705, 34.22798, 32.50315, 31.3762, 34.4286,
    36.57304, 32.63208, 32.20542, 33.74768, 33.67143, 31.2146, 28.97899,
    30.51925, 34.81638, 35.67587, 31.92131, 32.44133, 38.72983, 37.48034,
    28.37461, 26.34083,
  40.04165, 42.406, 44.14377, 45.93954, 45.32883, 41.21377, 36.63609,
    36.44854, 35.63729, 34.82164, 35.13963, 38.11618, 39.02428, 37.44145,
    35.01208, 34.96295, 35.71896, 36.15272, 34.63301, 32.8727, 33.03468,
    33.68692, 34.5997, 32.75113, 38.00229, 48.63285, 41.35519, 29.45756,
    26.77111, 25.49397,
  56.04807, 58.89183, 54.19416, 48.08484, 46.1208, 44.63268, 40.56473,
    42.21151, 43.7542, 51.2539, 55.91996, 39.35731, 34.25127, 33.17474,
    32.35479, 33.05209, 34.139, 34.06104, 32.92165, 32.74089, 35.30442,
    34.75261, 31.69895, 29.54818, 33.32686, 37.21297, 31.5762, 26.28456,
    25.87064, 25.32114,
  71.98257, 58.92411, 62.27565, 64.18007, 62.52682, 54.02674, 55.75024,
    52.0404, 43.99131, 47.73103, 46.84704, 33.29364, 33.89721, 34.54506,
    32.15955, 32.58031, 31.87334, 31.72358, 31.31386, 31.85571, 34.78939,
    33.5193, 29.11034, 32.57144, 34.62276, 28.26677, 25.79152, 26.15749,
    26.05828, 25.52442,
  80.79321, 79.00681, 89.24763, 91.90911, 94.19343, 89.92619, 68.56685,
    46.7742, 45.20966, 42.3046, 39.30064, 32.61748, 36.71648, 38.6546,
    33.73621, 32.57588, 32.43003, 31.83787, 30.93963, 33.12399, 34.824,
    31.56442, 28.6184, 33.42038, 34.94451, 27.37565, 26.01105, 26.30066,
    26.54235, 25.81134,
  87.43828, 92.59679, 93.56566, 93.02682, 84.16045, 74.55066, 73.59728,
    66.03102, 57.77373, 52.26875, 59.67744, 57.8423, 58.72936, 57.40812,
    49.8094, 39.67957, 33.05502, 34.6131, 35.86689, 36.88142, 33.89713,
    32.83714, 34.81643, 30.80272, 28.30663, 26.66769, 26.05938, 25.8608,
    26.24178, 25.77823,
  65.95442, 70.39769, 65.33325, 60.6132, 54.22313, 61.81144, 85.59699,
    82.65637, 72.2299, 73.25867, 69.76397, 53.88132, 43.01212, 47.99717,
    50.37669, 36.73042, 36.75102, 36.80751, 40.21115, 41.4438, 36.72493,
    33.31614, 30.08235, 27.43039, 26.39666, 26.75373, 26.15718, 25.7604,
    25.74964, 25.50655,
  52.51456, 50.64916, 49.04097, 47.22117, 47.34059, 52.62324, 59.27272,
    57.60383, 54.34095, 52.14608, 47.98165, 40.00875, 35.26955, 38.59463,
    38.55989, 35.93108, 37.44966, 35.93806, 37.19474, 36.97893, 31.25337,
    28.63501, 26.58775, 26.46344, 26.81115, 26.68232, 26.23719, 25.86843,
    25.68931, 25.42353,
  47.70678, 45.54974, 44.41015, 44.32625, 45.44365, 46.31213, 46.62465,
    46.45651, 44.92104, 42.29924, 37.55502, 36.4094, 39.88508, 38.40175,
    36.08897, 35.98331, 35.31801, 33.5518, 35.48239, 34.46592, 27.43479,
    27.47565, 27.10307, 26.62445, 26.56602, 26.67572, 26.17926, 25.64015,
    25.58867, 25.41805,
  43.36132, 43.04287, 42.69313, 43.26961, 43.42134, 43.74678, 43.55846,
    42.96218, 41.8093, 38.29251, 37.03071, 39.20123, 39.37819, 38.72345,
    40.01332, 37.53123, 33.15286, 30.6976, 33.83776, 32.95729, 27.53648,
    27.83375, 27.53422, 26.95844, 26.21177, 26.32125, 26.01717, 25.47055,
    25.42286, 25.33525,
  44.07169, 44.23108, 42.74901, 41.81094, 41.55612, 40.96798, 40.45713,
    39.89555, 38.32492, 36.3655, 37.83988, 37.7286, 33.53075, 33.99953,
    34.80565, 33.71436, 33.36317, 33.69109, 36.58212, 35.93676, 30.97578,
    28.80699, 27.76268, 27.16248, 26.14489, 25.98058, 25.82897, 25.47653,
    25.38349, 25.30492,
  44.5943, 44.19621, 42.18148, 40.26349, 39.74436, 39.20751, 38.74508,
    38.07675, 36.95157, 37.81731, 38.0358, 33.49935, 30.87102, 30.89882,
    30.65361, 30.00078, 31.40283, 33.51598, 35.75219, 36.74704, 34.21333,
    30.65091, 28.06917, 27.37313, 26.56095, 26.01527, 25.77382, 25.50607,
    25.38357, 25.31817,
  43.53808, 42.93085, 40.86908, 39.13924, 38.55379, 38.30338, 37.96728,
    37.28503, 36.79314, 37.52066, 34.83034, 30.07668, 30.03038, 30.32916,
    29.97499, 29.28308, 29.62575, 30.35327, 31.84213, 32.54106, 32.03555,
    31.40901, 29.88968, 28.08094, 26.93178, 26.27821, 25.7721, 25.50448,
    25.39776, 25.31577,
  43.38792, 41.68062, 39.98772, 38.82548, 38.32798, 37.63382, 37.26773,
    36.41396, 36.69341, 36.04121, 31.66181, 28.84768, 29.36645, 29.55955,
    29.39907, 29.16619, 28.82912, 28.75441, 29.00702, 28.81271, 29.95821,
    30.74525, 30.63017, 30.939, 29.00254, 26.82119, 25.8581, 25.63585,
    25.43596, 25.33062,
  42.31676, 41.15008, 39.2224, 38.11344, 38.47962, 38.53483, 37.76634,
    36.27453, 36.17068, 34.12447, 29.77988, 28.62192, 28.89391, 29.06184,
    28.788, 29.11253, 29.05033, 28.13887, 27.68702, 27.56073, 28.90153,
    29.32175, 28.57004, 30.20023, 30.40696, 27.83026, 26.12116, 26.09663,
    25.72325, 25.36479,
  41.47635, 40.49027, 39.60148, 39.11475, 39.0256, 38.74555, 38.81991,
    38.38459, 38.26606, 34.25843, 29.53457, 29.27016, 29.5621, 29.99533,
    29.88431, 29.85868, 30.04169, 29.18436, 27.93701, 27.77239, 28.19173,
    28.11469, 27.75243, 28.15998, 29.33698, 29.40761, 27.69537, 26.46642,
    26.08073, 25.51041,
  40.8978, 41.16048, 39.00126, 38.28964, 38.59839, 38.46416, 37.96601,
    37.9049, 38.77844, 34.83904, 29.73778, 29.62626, 30.08378, 30.35814,
    30.37137, 30.46355, 30.19892, 29.96129, 28.76794, 27.60114, 27.92582,
    28.19116, 28.01376, 27.38953, 27.11855, 28.43638, 28.57875, 27.25112,
    26.92309, 25.93828,
  40.86825, 42.51187, 41.65709, 39.8758, 38.62671, 37.7566, 38.73694,
    39.79676, 38.00107, 33.68289, 30.41231, 30.2652, 30.88919, 30.48852,
    29.82183, 29.88085, 29.77785, 29.82792, 29.06371, 27.83102, 28.32811,
    28.65149, 27.61847, 26.82368, 26.73987, 27.36424, 28.72473, 27.97621,
    26.81671, 25.82947,
  41.86309, 43.34155, 40.80183, 39.00441, 38.21315, 37.43232, 38.9246,
    39.42208, 35.85813, 32.11853, 30.65798, 30.53243, 30.68155, 30.1151,
    29.66598, 29.46904, 29.28312, 29.48972, 28.88934, 27.73048, 28.55981,
    30.14352, 30.18091, 28.86331, 28.29497, 28.47871, 30.20571, 29.95984,
    26.87917, 25.30799,
  41.39893, 41.52793, 39.62583, 39.04103, 39.4792, 39.19228, 39.76098,
    37.94939, 33.56764, 31.51452, 30.30823, 30.13799, 30.16319, 29.88856,
    30.10073, 29.83496, 29.18292, 29.22755, 29.32556, 29.23309, 30.72671,
    31.45829, 30.45702, 29.17537, 28.7312, 28.92836, 29.36534, 31.28129,
    29.71336, 26.08891,
  38.98964, 38.21818, 38.68906, 39.94258, 41.08716, 42.4044, 40.98806,
    36.56475, 33.12996, 31.5711, 29.55452, 28.5233, 28.40351, 29.01191,
    30.1151, 30.57795, 30.7248, 31.20292, 30.29628, 29.09785, 29.35707,
    29.01736, 27.96702, 27.3794, 27.59545, 28.09384, 28.21855, 28.2966,
    28.89235, 26.72271,
  38.02375, 38.22732, 38.33543, 38.22552, 38.75433, 41.53597, 42.10039,
    36.85569, 32.84751, 31.86402, 30.97486, 30.69419, 30.7774, 31.50867,
    32.19005, 32.21175, 31.19239, 29.86387, 28.91314, 27.78347, 27.19322,
    26.96678, 26.76657, 26.67448, 26.78523, 27.31435, 27.4374, 26.87999,
    26.41292, 25.58657,
  17.459, 17.49169, 17.52716, 17.54892, 17.5316, 17.52752, 17.53817,
    17.55175, 17.60316, 17.66378, 18.4222, 18.52825, 17.6692, 17.82196,
    17.94036, 17.64867, 17.57485, 17.60738, 17.61712, 18.08866, 18.34206,
    17.89672, 17.82693, 18.24978, 18.46403, 18.13296, 20.30568, 21.86584,
    19.23264, 18.10541,
  17.78685, 17.8265, 17.64215, 17.8749, 17.72684, 17.58619, 17.6365,
    17.68567, 17.76331, 17.90453, 18.25997, 18.75158, 19.03062, 18.43872,
    18.15072, 18.18997, 17.74025, 17.77371, 18.1611, 18.59336, 18.53592,
    18.02404, 18.00599, 18.60239, 22.24509, 23.04075, 21.03446, 24.21742,
    20.1895, 18.72223,
  17.72149, 17.73067, 17.69026, 17.74252, 17.69282, 17.65352, 17.66852,
    17.73236, 17.82638, 17.88613, 17.96892, 18.33939, 18.61533, 19.01733,
    19.11277, 18.36194, 18.264, 18.55927, 18.55937, 18.72991, 19.40283,
    20.55766, 21.46537, 20.94783, 25.65203, 28.72815, 23.5029, 23.93888,
    20.11771, 19.24282,
  17.72949, 17.72543, 17.88834, 18.03282, 18.24749, 18.67599, 18.72052,
    18.47849, 18.52648, 18.766, 18.84495, 19.13145, 18.96739, 18.65182,
    19.49127, 20.32329, 19.72094, 18.76196, 18.90334, 19.2265, 21.49031,
    22.8742, 21.90805, 26.16055, 28.17653, 25.30284, 26.35087, 23.43566,
    20.04162, 18.57172,
  18.19598, 17.95464, 18.19959, 18.51388, 18.80449, 18.97404, 18.9407,
    18.79734, 19.29302, 19.66865, 19.4485, 19.33938, 19.1717, 19.37464,
    20.00374, 20.48667, 19.72019, 19.0682, 19.48611, 23.89144, 25.65226,
    21.1431, 20.9986, 22.93793, 24.52048, 24.20542, 23.42094, 23.70187,
    24.25723, 20.13211,
  18.31715, 18.40729, 19.06351, 20.01254, 19.97177, 19.47676, 19.53209,
    19.35449, 19.05902, 19.14318, 19.14511, 20.7212, 22.70064, 22.83521,
    22.21547, 28.56238, 35.33947, 27.77125, 22.46848, 24.49882, 23.11417,
    19.91315, 20.33393, 21.14488, 23.67516, 23.40267, 25.54867, 37.16366,
    33.91994, 19.66379,
  18.84434, 19.16056, 19.8713, 20.7307, 20.81433, 20.51164, 21.19437,
    22.65018, 22.9288, 22.84473, 23.47666, 23.25418, 22.37872, 22.46895,
    27.17807, 34.3193, 32.26674, 24.86271, 22.35438, 22.08779, 20.70493,
    19.8515, 20.37578, 22.66762, 24.24469, 21.97652, 30.88352, 45.81245,
    34.28249, 18.21798,
  19.81866, 20.1897, 21.05514, 22.00388, 21.94641, 23.77729, 25.98486,
    24.24421, 22.79428, 22.87124, 22.76376, 21.89607, 20.97664, 21.16414,
    23.27233, 25.06577, 23.87094, 22.34634, 20.88164, 20.61794, 20.09608,
    19.83171, 21.1109, 23.45526, 23.29183, 21.71079, 34.11769, 40.13275,
    24.48998, 18.41205,
  22.52547, 22.81298, 23.88096, 24.23411, 24.63292, 26.40221, 25.61136,
    23.95411, 23.70741, 23.51003, 22.66306, 21.57127, 20.94901, 23.92501,
    25.8619, 22.71566, 22.5924, 24.133, 24.05372, 21.89017, 19.97065,
    21.32557, 25.31468, 26.16469, 22.908, 23.33889, 30.05489, 29.01937,
    20.39943, 18.44883,
  26.56787, 28.22883, 29.7554, 31.20553, 31.30413, 28.34022, 24.57619,
    24.21146, 23.45935, 22.51721, 23.00446, 25.94248, 27.41865, 27.04499,
    25.41865, 25.30653, 26.03018, 26.6037, 25.25745, 23.5498, 23.48022,
    24.28227, 25.48495, 24.07139, 28.81643, 38.2258, 32.06164, 21.46136,
    18.9333, 17.72352,
  38.93629, 42.32452, 39.03662, 34.35651, 33.02492, 31.61934, 27.89804,
    29.12362, 30.10712, 36.75577, 40.59324, 27.78481, 24.20886, 23.65135,
    22.93177, 23.74172, 24.9047, 24.91075, 23.77172, 23.43431, 25.74544,
    25.62349, 22.91854, 21.02872, 25.09168, 29.40404, 23.91782, 18.46947,
    18.03621, 17.55406,
  53.67579, 43.4983, 45.76135, 46.73243, 45.13575, 38.79174, 41.37333,
    38.60139, 31.59019, 35.88643, 35.58757, 22.77299, 23.50485, 24.26772,
    22.61251, 23.0462, 22.57669, 22.51497, 22.11112, 22.67817, 25.48338,
    24.53069, 20.65562, 23.79132, 25.73921, 20.36935, 17.99405, 18.29725,
    18.22197, 17.72627,
  61.64826, 57.7928, 74.70472, 79.76643, 80.62555, 71.84711, 55.31051,
    35.61943, 33.27384, 31.48523, 28.40946, 21.23547, 25.60128, 27.9707,
    23.86097, 23.07109, 23.1561, 22.53263, 21.92408, 24.10884, 25.85593,
    22.99617, 20.33459, 25.22264, 26.74267, 19.58801, 18.14238, 18.43369,
    18.67206, 17.98732,
  68.05116, 91.5593, 93.57806, 89.52888, 78.72385, 67.96196, 58.58939,
    51.92286, 43.74318, 38.18535, 43.65498, 42.01522, 44.69062, 44.3629,
    37.80016, 29.35897, 23.67846, 25.17744, 26.46972, 27.57113, 25.17432,
    24.1561, 25.91274, 23.08082, 20.59856, 18.73, 18.19586, 18.05471,
    18.44092, 17.97518,
  51.6348, 59.67702, 57.35268, 54.58045, 48.23885, 50.90853, 68.03174,
    66.24567, 56.37513, 56.49072, 54.71689, 41.97324, 32.91725, 38.07124,
    39.92651, 27.63158, 26.98711, 27.25507, 29.98832, 31.08227, 27.72097,
    25.04404, 22.44289, 19.77779, 18.40403, 18.76273, 18.27765, 17.94293,
    17.96683, 17.73147,
  40.7602, 40.40321, 39.50777, 37.68484, 36.61642, 40.74599, 47.51591,
    45.7365, 42.35234, 41.1531, 37.98632, 29.82114, 25.15134, 29.09993,
    29.15943, 26.49467, 28.07969, 26.72475, 27.70426, 27.66892, 23.29255,
    20.92465, 18.82089, 18.66569, 18.90761, 18.70063, 18.33397, 18.04098,
    17.90424, 17.65992,
  38.04622, 36.51679, 34.88992, 34.03424, 34.57753, 35.54372, 35.91577,
    35.61915, 34.20367, 31.79701, 27.17646, 26.11771, 29.26187, 27.83585,
    26.53845, 26.76798, 26.4623, 24.74184, 26.00514, 25.08569, 19.51181,
    19.44277, 19.19128, 18.84888, 18.7348, 18.7226, 18.27839, 17.85144,
    17.82693, 17.65834,
  34.16472, 33.16323, 32.20934, 32.59455, 32.97561, 33.69112, 33.86693,
    33.36768, 31.98617, 28.20017, 26.62535, 29.02168, 29.51443, 28.97523,
    30.40757, 28.55878, 24.76342, 22.48054, 24.9855, 23.99708, 19.44933,
    19.75644, 19.5731, 19.11896, 18.39204, 18.43875, 18.18318, 17.69874,
    17.67167, 17.58744,
  33.54288, 33.36642, 32.0623, 31.57492, 31.7618, 31.63903, 31.39956,
    30.70607, 28.75522, 26.4673, 27.99797, 28.39161, 24.93012, 25.59026,
    26.48382, 25.45256, 24.82233, 24.91496, 27.09572, 26.15614, 22.24946,
    20.64186, 19.76495, 19.24938, 18.29945, 18.14178, 18.02083, 17.70296,
    17.63149, 17.55832,
  33.85049, 33.78078, 32.18734, 30.7093, 30.58939, 30.27533, 29.82507,
    29.0496, 27.78074, 28.49617, 29.00186, 25.21272, 22.71895, 22.75034,
    22.49046, 21.84173, 22.95306, 24.81321, 26.48151, 27.04467, 25.30134,
    22.40139, 19.97634, 19.3729, 18.64332, 18.16989, 17.97605, 17.73377,
    17.62894, 17.5622,
  33.34805, 33.33096, 31.60708, 30.09018, 29.72116, 29.60629, 29.37456,
    28.84677, 28.49785, 29.41528, 27.08682, 22.38845, 22.06024, 22.06328,
    21.51051, 20.84949, 21.1885, 21.99937, 23.18979, 23.77394, 23.72273,
    23.19945, 21.61628, 19.99785, 18.99207, 18.40129, 17.96365, 17.73375,
    17.64762, 17.56645,
  33.73626, 32.66413, 31.08859, 30.09595, 29.81884, 29.43633, 29.48554,
    29.05767, 29.35862, 28.74424, 24.37, 21.05061, 21.22767, 21.20233,
    20.92746, 20.76241, 20.55245, 20.53203, 20.86698, 20.79276, 21.83235,
    22.28028, 21.79586, 22.10925, 20.68682, 18.84654, 18.05867, 17.83626,
    17.67396, 17.57472,
  33.34002, 32.52248, 30.7436, 29.88039, 30.52187, 30.96446, 30.73138,
    29.5582, 29.29752, 27.05475, 22.39733, 20.63617, 20.6153, 20.6762,
    20.44344, 20.81989, 20.7913, 20.00653, 19.67774, 19.58196, 20.81178,
    20.93487, 20.00384, 21.65124, 21.99482, 19.7111, 18.29046, 18.23912,
    17.9153, 17.59961,
  32.86579, 32.22595, 31.46912, 31.35197, 31.73011, 31.87365, 32.04807,
    31.41779, 30.87756, 26.76995, 21.88485, 21.12923, 21.22588, 21.56962,
    21.44917, 21.51142, 21.63331, 20.7843, 19.79103, 19.7335, 20.07899,
    19.8945, 19.46685, 19.91366, 21.06378, 21.16722, 19.69934, 18.59276,
    18.24905, 17.72207,
  32.87598, 33.67009, 31.72899, 31.2267, 31.68793, 31.57009, 31.0667,
    30.80319, 31.30631, 27.22905, 22.10828, 21.54276, 21.6917, 21.96234,
    22.00843, 22.04094, 21.68106, 21.29162, 20.40432, 19.6253, 19.76068,
    19.8512, 19.73066, 19.24922, 19.16675, 20.43338, 20.54845, 19.30144,
    19.045, 18.11329,
  33.41739, 35.54973, 34.1844, 32.52779, 31.44743, 30.55136, 31.21216,
    32.09865, 30.64442, 26.38808, 22.79432, 22.13053, 22.34913, 22.03628,
    21.50392, 21.52217, 21.24157, 21.11819, 20.65847, 19.79776, 20.05966,
    20.23568, 19.43834, 18.8304, 18.77991, 19.39551, 20.68466, 19.94238,
    19.00569, 18.04469,
  34.47039, 36.35873, 33.73923, 31.7515, 30.79807, 29.90057, 31.37605,
    32.09816, 28.89708, 25.03462, 23.13748, 22.44266, 22.22221, 21.70493,
    21.28024, 21.09534, 20.83707, 20.86466, 20.51212, 19.70944, 20.151,
    21.29249, 21.27776, 20.40345, 20.18838, 20.34894, 22.06578, 21.73086,
    18.98884, 17.59556,
  34.03313, 34.4839, 32.25425, 31.31718, 31.65031, 31.30789, 32.11197,
    30.84507, 26.8783, 24.46932, 22.82886, 22.05416, 21.70262, 21.47418,
    21.7093, 21.44095, 20.73428, 20.59408, 20.83336, 20.99446, 21.80411,
    22.12644, 21.53537, 20.76461, 20.69175, 20.81123, 21.32202, 23.09748,
    21.50455, 18.21807,
  31.47744, 30.69702, 30.98587, 32.18007, 33.24773, 34.33415, 33.35585,
    29.6024, 26.30176, 24.42482, 22.04599, 20.61524, 20.27395, 20.61646,
    21.41067, 21.71753, 21.6761, 22.01446, 21.57322, 20.92638, 21.05754,
    20.7071, 19.85055, 19.40149, 19.64708, 20.10517, 20.19728, 20.3807,
    20.96852, 18.77814,
  30.10525, 30.30711, 30.59955, 30.78301, 31.29275, 33.69395, 34.11783,
    29.50173, 25.78126, 24.35157, 22.88663, 22.17262, 22.16316, 22.51543,
    22.84668, 22.9335, 22.13812, 21.15151, 20.54627, 19.74851, 19.24779,
    19.11118, 18.9084, 18.78831, 18.88454, 19.40146, 19.54327, 19.00219,
    18.62468, 17.83346,
  11.62529, 11.65557, 11.6851, 11.70018, 11.68632, 11.68294, 11.69184,
    11.70097, 11.73932, 11.76237, 12.4777, 12.54015, 11.78791, 11.95212,
    12.05672, 11.79388, 11.71955, 11.7434, 11.74752, 12.18207, 12.40316,
    12.02786, 11.97063, 12.32057, 12.43393, 12.08506, 14.2093, 15.62098,
    13.38862, 12.24155,
  11.92103, 11.93445, 11.80216, 12.00084, 11.85759, 11.73069, 11.7617,
    11.80179, 11.86137, 11.98444, 12.35873, 12.81491, 13.02172, 12.49059,
    12.28586, 12.27428, 11.85918, 11.87541, 12.23249, 12.64536, 12.58936,
    12.05939, 11.98994, 12.48374, 15.83603, 16.32878, 15.17103, 18.01794,
    14.32131, 12.83309,
  11.87512, 11.87466, 11.83799, 11.88544, 11.81803, 11.75386, 11.76246,
    11.81938, 11.90032, 11.95884, 12.03023, 12.39329, 12.68056, 13.04613,
    13.07649, 12.36283, 12.27779, 12.53223, 12.49052, 12.57672, 13.09234,
    14.07646, 14.87265, 14.26305, 18.94036, 21.69124, 17.28108, 17.75427,
    14.16106, 13.28965,
  11.83397, 11.8162, 11.95621, 12.07097, 12.25883, 12.62459, 12.64729,
    12.42605, 12.45043, 12.67829, 12.76569, 13.02722, 12.81052, 12.59641,
    13.36097, 14.06263, 13.47358, 12.54955, 12.50389, 12.60497, 14.74423,
    16.03912, 15.27147, 19.17911, 20.94591, 19.00199, 20.02639, 17.31532,
    14.04487, 12.66847,
  12.17958, 11.92672, 12.13464, 12.42024, 12.71494, 12.86016, 12.78294,
    12.61705, 13.13314, 13.6089, 13.49734, 13.24167, 12.90349, 13.05438,
    13.67334, 14.00848, 13.06229, 12.37287, 12.64927, 16.86083, 18.4107,
    14.49973, 14.4313, 16.54061, 18.03249, 17.65725, 17.1018, 17.44025,
    17.66407, 13.8529,
  12.12119, 12.11897, 12.75735, 13.73738, 13.7904, 13.26562, 13.17036,
    12.96525, 12.75511, 12.87908, 12.7865, 14.12972, 15.74629, 15.88449,
    15.1235, 20.92189, 26.70972, 19.88025, 15.29738, 17.64294, 16.43509,
    13.40243, 13.9184, 14.55056, 16.903, 16.5041, 18.76934, 29.83244,
    26.54791, 13.46781,
  12.17512, 12.44735, 13.22206, 14.1626, 14.3437, 13.8843, 14.29113,
    15.65408, 15.92735, 15.82173, 16.42282, 16.18677, 15.35871, 15.24198,
    19.79626, 26.79988, 24.94884, 17.78157, 15.55008, 15.45331, 14.20731,
    13.40919, 13.82392, 15.7922, 17.26304, 14.9859, 23.63969, 38.1816,
    27.42103, 12.21666,
  12.34696, 12.65986, 13.55159, 14.42524, 14.33418, 16.06638, 17.9831,
    16.39738, 15.2683, 15.47897, 15.58643, 14.70604, 13.74747, 13.87068,
    16.43039, 18.49052, 17.04152, 15.46451, 14.35495, 14.13821, 13.66266,
    13.40001, 14.41614, 16.54658, 16.50279, 14.57893, 27.1499, 33.33961,
    18.18802, 12.41632,
  13.7353, 13.86186, 14.92429, 15.14447, 15.57551, 17.55635, 16.93795,
    15.25113, 15.29713, 15.53476, 15.01263, 14.1041, 13.6397, 16.63629,
    18.39757, 15.69773, 15.62815, 16.93909, 16.86266, 15.00735, 13.37264,
    14.41795, 17.91412, 18.84612, 16.07395, 15.99669, 22.74986, 22.28598,
    14.10848, 12.49793,
  15.88534, 17.10299, 18.65457, 19.99244, 20.39281, 17.91495, 14.76172,
    14.58061, 14.4168, 13.88158, 14.87518, 17.93747, 19.27776, 19.213,
    18.30529, 18.1044, 18.65028, 19.14536, 18.30448, 17.06747, 16.8613,
    17.71858, 19.04246, 17.75219, 21.81267, 30.32367, 25.00446, 15.41478,
    13.05054, 11.86862,
  25.25292, 28.23217, 25.87579, 21.83983, 21.04239, 20.19479, 17.34578,
    18.88025, 20.28051, 26.5839, 29.88263, 19.86922, 17.16213, 16.75166,
    16.18646, 17.07605, 18.31002, 18.41564, 17.45724, 17.32755, 19.55242,
    19.57783, 17.05193, 15.10048, 19.11103, 23.74116, 18.50591, 12.75352,
    12.1641, 11.69464,
  38.42037, 29.42782, 30.8635, 31.63739, 30.2662, 26.15366, 29.17589,
    27.15585, 21.98095, 26.76752, 26.81337, 15.81288, 16.62162, 17.55481,
    16.28301, 16.74248, 16.39128, 16.39689, 16.09824, 16.68942, 19.46304,
    18.58834, 14.74217, 17.71808, 19.82423, 14.71817, 12.18532, 12.39868,
    12.32672, 11.8573,
  44.24705, 40.89961, 57.93153, 63.07863, 63.06326, 55.09444, 41.01857,
    25.80339, 23.96008, 23.14401, 20.24452, 14.2087, 18.77957, 21.1354,
    17.50363, 16.86565, 16.95699, 16.35405, 15.85314, 18.16797, 19.94879,
    17.02449, 14.34835, 19.46083, 21.24393, 13.82351, 12.2465, 12.5528,
    12.79098, 12.13813,
  53.14084, 77.37314, 78.26319, 73.0516, 62.22615, 53.41011, 47.15095,
    40.57726, 33.02, 28.45593, 33.36687, 32.70535, 36.0707, 36.08859,
    30.32225, 22.7288, 17.40705, 18.78046, 20.07837, 21.29028, 19.09364,
    18.11845, 19.92854, 17.48684, 15.03492, 12.8399, 12.3238, 12.19514,
    12.58208, 12.13814,
  39.80044, 48.41353, 46.48499, 43.56897, 37.19534, 40.5051, 56.16457,
    54.06133, 45.0481, 44.95261, 44.84448, 34.18109, 26.01387, 31.11128,
    33.19725, 21.29666, 20.42062, 20.50573, 22.3622, 23.84988, 21.85948,
    19.32141, 17.04047, 14.19108, 12.4377, 12.81076, 12.38947, 12.08288,
    12.11319, 11.88744,
  28.99938, 29.11711, 28.99737, 28.00414, 27.09245, 31.74125, 38.93361,
    36.75733, 33.97071, 33.92031, 31.02736, 23.44666, 18.60433, 22.75912,
    23.02002, 19.99413, 21.63018, 20.04091, 20.30559, 20.72077, 17.67717,
    15.41803, 13.1792, 12.99838, 13.06405, 12.75526, 12.42075, 12.17586,
    12.04397, 11.81065,
  27.08603, 26.358, 25.21835, 24.46225, 24.84661, 25.91636, 26.71627,
    26.51652, 25.92586, 24.70511, 20.66862, 19.94617, 22.30284, 20.7468,
    20.11599, 20.39684, 20.25911, 18.31791, 18.90379, 18.29727, 13.6479,
    13.5925, 13.41426, 13.20189, 12.95791, 12.78229, 12.36757, 11.99598,
    11.9634, 11.80243,
  24.36067, 23.61805, 22.60637, 22.84108, 23.31212, 24.23747, 24.92561,
    25.11567, 24.47314, 21.72398, 20.28424, 22.63811, 23.2596, 22.34833,
    23.93913, 22.38515, 18.79588, 16.38482, 18.32147, 17.42281, 13.46997,
    13.72567, 13.61501, 13.31939, 12.58506, 12.53489, 12.29616, 11.83847,
    11.80966, 11.72702,
  23.94803, 23.77312, 22.45885, 22.1423, 22.58292, 22.94658, 23.2955,
    23.21107, 21.94509, 20.21913, 21.70386, 22.33032, 19.26318, 19.80497,
    20.75114, 19.72306, 18.83184, 18.60682, 20.08897, 18.97169, 15.83878,
    14.54092, 13.69459, 13.30194, 12.4303, 12.25421, 12.15407, 11.83561,
    11.76567, 11.7022,
  24.28332, 24.338, 22.94098, 21.80315, 22.02637, 22.04521, 21.99751,
    21.72474, 20.91662, 21.89732, 22.82535, 19.59439, 17.12848, 17.01667,
    16.73076, 16.2086, 17.12107, 18.69094, 19.56932, 19.71567, 18.68494,
    16.24213, 13.8437, 13.4099, 12.75012, 12.2846, 12.10368, 11.86732,
    11.76943, 11.7078,
  23.94528, 24.26097, 22.9048, 21.70259, 21.56119, 21.55964, 21.47488,
    21.32602, 21.46128, 23.01512, 21.56103, 17.15759, 16.68863, 16.32315,
    15.52334, 14.9211, 15.20727, 15.96842, 16.65205, 16.99514, 17.4722,
    17.18608, 15.40405, 14.01674, 13.14344, 12.5321, 12.10481, 11.86581,
    11.77371, 11.70848,
  24.55725, 24.08848, 22.77461, 21.95959, 21.72107, 21.28952, 21.46119,
    21.50691, 22.39426, 22.84535, 19.4302, 15.89976, 15.75062, 15.37975,
    14.86846, 14.67307, 14.48672, 14.44593, 14.78724, 14.7898, 15.92982,
    16.27315, 15.3758, 15.6682, 14.50418, 12.89796, 12.1861, 11.95409,
    11.7887, 11.71154,
  24.66828, 24.27429, 22.61007, 21.75889, 22.2604, 22.61798, 22.73689,
    22.18586, 22.64999, 21.56997, 17.55783, 15.38472, 14.97287, 14.72991,
    14.36811, 14.70543, 14.68464, 13.99124, 13.79743, 13.76534, 15.01564,
    14.95256, 13.70399, 15.28339, 15.65527, 13.66079, 12.41591, 12.35428,
    12.03318, 11.73257,
  24.40733, 24.07138, 23.16238, 22.99055, 23.48823, 23.81981, 24.43435,
    24.33122, 24.25573, 21.05841, 16.77567, 15.67256, 15.39579, 15.44924,
    15.1775, 15.29326, 15.42318, 14.62473, 13.83509, 13.8908, 14.17604,
    13.8439, 13.33327, 13.74802, 14.77, 15.04499, 13.79403, 12.70967,
    12.37477, 11.85954,
  24.55334, 25.27538, 23.44543, 23.06731, 23.82376, 24.02942, 23.84562,
    23.78557, 24.49847, 21.27769, 16.76827, 15.92539, 15.66662, 15.78251,
    15.79651, 15.81178, 15.43332, 14.99993, 14.32809, 13.82243, 13.76547,
    13.69726, 13.63792, 13.2495, 13.23492, 14.5644, 14.71882, 13.45092,
    13.19186, 12.26367,
  25.04421, 27.17619, 25.85289, 24.3909, 23.90599, 23.27234, 23.72345,
    24.55079, 23.616, 20.42644, 17.31256, 16.39993, 16.20456, 15.86678,
    15.37612, 15.32732, 14.96955, 14.79276, 14.55504, 13.94356, 13.97367,
    14.04016, 13.4133, 12.91701, 12.90774, 13.55903, 14.8564, 14.09764,
    13.21693, 12.27105,
  26.24703, 28.56019, 26.22442, 24.20689, 23.32143, 22.33864, 23.80488,
    24.66324, 22.07165, 19.1338, 17.73722, 16.82183, 16.19467, 15.58459,
    15.07493, 14.85816, 14.58604, 14.57298, 14.4251, 13.85869, 14.01749,
    14.8784, 14.89544, 14.33379, 14.28402, 14.45768, 16.23966, 15.86751,
    13.17671, 11.81085,
  26.48425, 27.50428, 24.94403, 23.5302, 23.64556, 23.0818, 23.9842,
    23.37633, 20.34398, 18.70234, 17.57178, 16.47957, 15.60577, 15.25616,
    15.40779, 15.13572, 14.47669, 14.29615, 14.70689, 15.09997, 15.4637,
    15.52852, 15.1489, 14.72041, 14.87471, 14.97991, 15.573, 17.32199,
    15.68552, 12.3858,
  24.4493, 23.5379, 23.42262, 24.48243, 25.18046, 25.58218, 24.92431,
    22.14583, 19.7424, 18.63605, 16.66217, 15.05984, 14.44189, 14.50452,
    15.05213, 15.26766, 15.17438, 15.44855, 15.34258, 15.04468, 15.05151,
    14.66411, 13.89398, 13.52001, 13.8199, 14.30088, 14.42932, 14.68847,
    15.22085, 12.95876,
  22.88921, 22.72359, 23.02512, 23.4687, 23.86234, 25.54858, 25.60361,
    21.95836, 19.19236, 18.32963, 17.00958, 16.23282, 16.18164, 16.11327,
    16.11261, 16.25491, 15.60286, 14.81323, 14.46016, 13.83623, 13.3743,
    13.28127, 13.06097, 12.93476, 13.04169, 13.57463, 13.78723, 13.22573,
    12.80195, 12.0114,
  10.94995, 10.97038, 11.00348, 11.01271, 11.00065, 11.00156, 11.00248,
    11.00786, 11.04206, 11.05127, 11.70676, 11.78197, 11.0768, 11.22859,
    11.33839, 11.09849, 11.0368, 11.05336, 11.03806, 11.42947, 11.65087,
    11.31286, 11.247, 11.5663, 11.6284, 11.2632, 13.23231, 14.55785,
    12.59402, 11.56276,
  11.21595, 11.22603, 11.10118, 11.30132, 11.16952, 11.04462, 11.07323,
    11.09514, 11.14932, 11.26148, 11.66963, 12.10159, 12.23397, 11.75219,
    11.56462, 11.55279, 11.15347, 11.15429, 11.48319, 11.93277, 11.90208,
    11.34553, 11.23052, 11.6855, 14.69019, 15.04816, 14.53333, 17.43943,
    13.68948, 12.18842,
  11.20881, 11.2062, 11.1501, 11.21856, 11.134, 11.04895, 11.05068, 11.10973,
    11.19954, 11.26025, 11.31882, 11.68145, 11.99406, 12.2791, 12.28979,
    11.62089, 11.50767, 11.76573, 11.75481, 11.82061, 12.20648, 13.03227,
    13.78043, 13.14757, 17.6481, 20.43294, 16.60906, 17.27846, 13.53342,
    12.66356,
  11.14202, 11.11802, 11.24388, 11.32919, 11.48786, 11.83403, 11.86207,
    11.65381, 11.66656, 11.87249, 11.9561, 12.23021, 12.02634, 11.83731,
    12.55193, 13.17318, 12.65706, 11.78483, 11.65392, 11.59769, 13.58649,
    14.94694, 14.24061, 17.94965, 19.83471, 18.33093, 19.50649, 16.77399,
    13.40158, 12.05761,
  11.4521, 11.19194, 11.36913, 11.61967, 11.91799, 12.0975, 12.02773,
    11.83542, 12.31133, 12.83711, 12.79726, 12.48604, 12.07726, 12.183,
    12.81997, 13.16286, 12.09843, 11.34051, 11.5361, 15.48355, 17.17968,
    13.64311, 13.49396, 15.8182, 17.30848, 16.79467, 16.55704, 16.79324,
    16.82708, 13.09402,
  11.38347, 11.31641, 11.89119, 12.81081, 12.95763, 12.48431, 12.34169,
    12.15495, 11.99027, 12.13404, 11.98001, 13.13361, 14.6152, 14.75264,
    13.86251, 18.89937, 24.23449, 18.20664, 14.00851, 16.62261, 15.67754,
    12.57654, 13.12909, 13.71185, 15.99554, 15.70796, 17.15483, 27.62037,
    25.47952, 12.84217,
  11.36548, 11.60577, 12.35283, 13.29249, 13.55433, 13.03947, 13.2462,
    14.52749, 14.74195, 14.60053, 15.15713, 15.04211, 14.3384, 14.0704,
    18.17661, 25.28931, 24.0667, 16.88656, 14.64479, 14.65497, 13.42869,
    12.64718, 13.0378, 14.88773, 16.39329, 14.04188, 22.10024, 37.23447,
    27.34149, 11.55385,
  11.4953, 11.7911, 12.63118, 13.46509, 13.34173, 14.83129, 16.63761,
    15.32588, 14.3034, 14.48043, 14.65189, 13.73684, 12.64874, 12.63409,
    15.42095, 17.91411, 16.32446, 14.53337, 13.56613, 13.40567, 12.95074,
    12.66019, 13.56699, 15.65334, 15.70046, 13.51138, 26.45525, 33.76532,
    17.88214, 11.71535,
  12.61545, 12.69686, 13.67517, 13.85057, 14.17949, 16.35368, 15.98237,
    14.12711, 14.12722, 14.38828, 13.86317, 12.89142, 12.3653, 15.29833,
    17.16431, 14.69344, 14.72128, 16.05117, 15.94786, 14.21587, 12.59487,
    13.48762, 16.82689, 17.86548, 15.17402, 14.89138, 22.15036, 22.13676,
    13.28363, 11.8504,
  14.21882, 15.23425, 16.81027, 18.19917, 18.64739, 16.44299, 13.45229,
    13.189, 13.13128, 12.58361, 13.43229, 16.38988, 17.81998, 18.04759,
    17.36309, 17.02895, 17.51462, 18.08804, 17.47684, 16.32001, 15.95795,
    16.83924, 18.30339, 17.07951, 20.57716, 28.92315, 24.39405, 14.91048,
    12.46437, 11.21791,
  21.68476, 24.56182, 22.94055, 19.38094, 18.91444, 18.09092, 15.31181,
    16.75581, 17.89163, 23.68224, 27.14815, 18.66072, 16.39919, 15.99789,
    15.35782, 16.25974, 17.52344, 17.63461, 16.70382, 16.60201, 18.81882,
    18.93815, 16.46922, 14.42388, 18.50517, 23.61109, 18.51126, 12.23122,
    11.52833, 11.01922,
  33.04828, 25.30704, 26.37515, 26.61257, 25.32925, 21.71523, 24.86873,
    23.6417, 19.33476, 24.44773, 25.18018, 14.92206, 15.59659, 16.60839,
    15.53569, 16.00725, 15.66407, 15.65635, 15.3474, 15.96283, 18.85353,
    18.0507, 14.09058, 16.96624, 19.39688, 14.43694, 11.61907, 11.72411,
    11.65853, 11.18812,
  42.0141, 35.41802, 45.08094, 50.5941, 50.96482, 45.54702, 34.65675,
    21.88425, 20.7901, 20.66934, 18.27743, 13.11193, 17.59469, 20.03142,
    16.7364, 16.06348, 16.1838, 15.56656, 15.11104, 17.56714, 19.51132,
    16.48662, 13.72381, 19.06294, 21.18251, 13.35229, 11.56989, 11.88031,
    12.12474, 11.4883,
  47.69605, 67.25895, 68.68269, 69.10497, 65.02571, 54.59698, 39.07183,
    34.91697, 27.61034, 23.88356, 29.06288, 29.58379, 33.26864, 33.79874,
    28.92682, 21.93903, 16.66112, 18.08618, 19.49221, 20.8575, 18.69444,
    17.64636, 19.73512, 17.40769, 14.74949, 12.1938, 11.65226, 11.53566,
    11.93397, 11.50027,
  32.85123, 41.25909, 41.8259, 42.47135, 38.26841, 38.40871, 49.57431,
    48.82798, 38.00357, 38.487, 39.87365, 31.31719, 24.7671, 29.70272,
    32.03104, 20.6402, 19.75849, 19.81127, 21.47701, 23.1462, 21.37245,
    19.1108, 17.06329, 13.89598, 11.73324, 12.12825, 11.72984, 11.41937,
    11.44774, 11.23621,
  22.11701, 22.61753, 23.53152, 23.13504, 21.47817, 25.66796, 33.6377,
    31.05014, 28.1475, 29.62388, 28.25719, 21.73405, 17.60901, 21.99081,
    22.31756, 19.35975, 21.13289, 19.43038, 19.44776, 20.15492, 17.42058,
    15.17077, 12.68794, 12.38182, 12.4229, 12.09974, 11.75949, 11.53033,
    11.3789, 11.14188,
  20.67454, 20.24496, 19.4721, 18.60515, 18.5332, 19.58931, 20.50329,
    20.18564, 20.51307, 20.83801, 18.1398, 18.27112, 21.04894, 19.78107,
    19.52879, 19.88612, 19.88733, 17.83782, 18.24829, 17.86335, 13.21507,
    13.03971, 12.79525, 12.63034, 12.36126, 12.14642, 11.71282, 11.34395,
    11.30149, 11.13585,
  18.39345, 17.72916, 16.72749, 16.81718, 17.24048, 18.11933, 18.89938,
    19.3834, 19.24179, 17.61299, 17.16451, 20.60834, 22.31903, 21.63863,
    23.52734, 22.07515, 18.47357, 15.84023, 17.67597, 16.93075, 12.81384,
    12.98569, 12.91983, 12.71451, 11.9887, 11.89573, 11.64939, 11.17091,
    11.14326, 11.06247,
  18.12811, 17.82232, 16.41312, 16.00627, 16.4765, 16.94707, 17.37561,
    17.43365, 16.61139, 15.82352, 18.4275, 20.45121, 18.51815, 19.41173,
    20.57187, 19.52044, 18.40341, 17.74548, 19.16963, 18.11302, 14.98993,
    13.78865, 12.96078, 12.64237, 11.78269, 11.58739, 11.49852, 11.16791,
    11.09351, 11.03054,
  18.45375, 18.30295, 16.85315, 15.70371, 15.95311, 15.98711, 15.94341,
    15.75658, 15.40306, 17.36478, 19.71333, 17.98184, 16.37745, 16.58915,
    16.4106, 15.91672, 16.69241, 17.9568, 18.62446, 18.89385, 17.93668,
    15.54029, 13.09247, 12.69597, 12.08425, 11.60777, 11.43088, 11.19904,
    11.09372, 11.03272,
  17.98178, 18.11499, 16.8117, 15.61976, 15.49886, 15.44328, 15.28156,
    15.24148, 15.93952, 18.66451, 18.79612, 15.75584, 16.03233, 15.89688,
    15.07225, 14.43342, 14.60035, 15.23586, 15.86513, 16.37822, 17.02568,
    16.55003, 14.46586, 13.2872, 12.50945, 11.86713, 11.44109, 11.19797,
    11.09808, 11.03702,
  18.52654, 17.89157, 16.61573, 15.80067, 15.5656, 15.07064, 15.20904,
    15.51224, 17.07553, 18.84517, 17.00631, 14.54197, 15.06158, 14.8885,
    14.32255, 14.01469, 13.78809, 13.772, 14.20881, 14.281, 15.409, 15.67849,
    14.57495, 14.87108, 13.74432, 12.20413, 11.49749, 11.27693, 11.11158,
    11.03084,
  18.63754, 17.99565, 16.39132, 15.53889, 15.99584, 16.30738, 16.5739,
    16.39928, 17.54699, 17.7977, 15.22974, 13.98152, 14.16433, 14.10828,
    13.72725, 13.99369, 14.01087, 13.38268, 13.23635, 13.23854, 14.44257,
    14.3445, 13.01036, 14.51422, 14.8344, 12.93078, 11.70162, 11.65449,
    11.35621, 11.06009,
  18.35687, 17.84132, 16.85896, 16.62233, 17.22214, 17.69601, 18.59188,
    18.93399, 19.35347, 17.16345, 14.26027, 14.13663, 14.40928, 14.69819,
    14.45186, 14.54735, 14.70117, 13.93131, 13.15008, 13.25435, 13.55946,
    13.17812, 12.60172, 12.98911, 13.97081, 14.22472, 13.02665, 12.01771,
    11.70149, 11.18496,
  18.33739, 18.56385, 17.08478, 16.90588, 17.88725, 18.44934, 18.52334,
    18.57245, 19.48661, 17.24893, 14.06213, 14.30589, 14.69859, 15.04062,
    15.04535, 15.04188, 14.70748, 14.27768, 13.63076, 13.1995, 13.09167,
    12.96291, 12.92774, 12.54989, 12.53714, 13.89854, 14.07331, 12.78943,
    12.52092, 11.61369,
  18.68717, 20.15468, 19.31099, 18.38001, 18.33047, 18.11409, 18.55944,
    19.28646, 18.44098, 16.32195, 14.45149, 14.70446, 15.20525, 15.11725,
    14.63196, 14.57296, 14.2284, 14.06453, 13.87797, 13.31285, 13.28456,
    13.32185, 12.72974, 12.24486, 12.22839, 12.91737, 14.23759, 13.47588,
    12.58309, 11.64587,
  19.91787, 21.73282, 20.13603, 18.65812, 17.94382, 17.17372, 18.81356,
    19.54492, 16.93544, 14.98563, 14.85964, 15.16289, 15.28891, 14.87393,
    14.31694, 14.06469, 13.83368, 13.86598, 13.76523, 13.2181, 13.31153,
    14.12179, 14.15094, 13.61596, 13.59001, 13.78893, 15.61409, 15.26895,
    12.53844, 11.16411,
  20.68814, 21.58078, 19.21072, 18.06709, 18.184, 17.68124, 18.5915, 17.8888,
    15.10912, 14.50086, 14.82092, 14.98807, 14.7814, 14.51828, 14.58652,
    14.32386, 13.72632, 13.57143, 13.99675, 14.41494, 14.71345, 14.79208,
    14.46364, 14.07773, 14.25676, 14.37079, 15.03312, 16.7907, 15.08446,
    11.72647,
  19.27605, 18.30963, 18.11791, 19.25889, 19.63628, 19.55935, 18.93065,
    16.33188, 14.47078, 14.53756, 14.08807, 13.71071, 13.63007, 13.77748,
    14.29649, 14.4931, 14.38864, 14.66077, 14.65131, 14.43591, 14.43242,
    14.03994, 13.26897, 12.89987, 13.22044, 13.70709, 13.84508, 14.1975,
    14.73594, 12.37382,
  18.17926, 17.78631, 18.099, 18.61496, 18.71059, 19.81959, 19.65778,
    16.34386, 14.27693, 14.55893, 14.54085, 14.7426, 15.13948, 15.21913,
    15.26133, 15.41235, 14.84158, 14.13251, 13.82272, 13.22331, 12.76146,
    12.6696, 12.43871, 12.29145, 12.40899, 12.96411, 13.19946, 12.6295,
    12.23084, 11.39585,
  10.61548, 10.63374, 10.66829, 10.67774, 10.66817, 10.66475, 10.66721,
    10.67542, 10.70232, 10.70209, 11.34921, 11.4332, 10.73468, 10.88941,
    11.0006, 10.7694, 10.7146, 10.7212, 10.69053, 11.07474, 11.31147,
    10.9823, 10.91687, 11.23207, 11.27176, 10.86211, 12.85231, 14.24101,
    12.29256, 11.28225,
  10.87461, 10.88557, 10.76278, 10.96751, 10.8413, 10.7156, 10.73585,
    10.75574, 10.80786, 10.91485, 11.41165, 11.855, 11.91065, 11.45174,
    11.2718, 11.24717, 10.82909, 10.80917, 11.14226, 11.65049, 11.66582,
    11.0562, 10.87632, 11.31123, 14.27264, 14.64885, 14.44455, 17.68545,
    13.62056, 11.99191,
  10.8988, 10.89698, 10.83032, 10.92283, 10.82133, 10.71536, 10.70914,
    10.76784, 10.86458, 10.94878, 11.01327, 11.41348, 11.7963, 12.03312,
    12.00105, 11.31202, 11.16257, 11.44478, 11.47475, 11.55186, 11.85653,
    12.59441, 13.3132, 12.53647, 17.42364, 20.74947, 16.66674, 17.63468,
    13.46131, 12.5088,
  10.81153, 10.78554, 10.91887, 10.99348, 11.13281, 11.48186, 11.50907,
    11.30567, 11.31622, 11.51333, 11.62733, 11.94394, 11.72703, 11.5657,
    12.29389, 12.86117, 12.38043, 11.53288, 11.32543, 11.14239, 13.10951,
    14.56899, 13.79974, 17.70433, 20.08819, 18.6402, 19.90969, 17.04278,
    13.30377, 11.87563,
  11.13625, 10.86195, 11.02687, 11.26408, 11.57118, 11.82056, 11.74557,
    11.49558, 11.97702, 12.5786, 12.59317, 12.25635, 11.76013, 11.82579,
    12.56502, 13.02426, 11.8397, 10.88647, 11.00361, 14.82658, 16.71341,
    13.32721, 13.03848, 15.83005, 17.54015, 16.82745, 16.82812, 16.88646,
    16.77139, 12.87074,
  11.07563, 10.93527, 11.48987, 12.42114, 12.6424, 12.19383, 12.01187,
    11.82222, 11.72766, 11.92295, 11.70886, 12.76111, 14.22855, 14.42548,
    13.55436, 18.05009, 23.10828, 17.52471, 13.40096, 16.34567, 15.53592,
    12.16103, 12.79274, 13.44444, 15.94232, 15.78424, 16.7488, 27.4585,
    25.90057, 12.72873,
  10.9739, 11.18369, 11.98296, 13.02534, 13.35895, 12.77151, 12.85118,
    14.10866, 14.27504, 14.09707, 14.62486, 14.6825, 14.15398, 13.81176,
    17.53504, 24.76949, 24.19588, 16.79673, 14.31434, 14.43241, 13.13442,
    12.29426, 12.76118, 14.74968, 16.44191, 13.86692, 21.90174, 38.4672,
    28.80797, 11.35204,
  11.09191, 11.39269, 12.29909, 13.19295, 13.0379, 14.40088, 16.24683,
    15.07561, 14.04374, 14.22693, 14.50003, 13.5331, 12.24958, 12.08161,
    15.12475, 18.04618, 16.31343, 14.20209, 13.24121, 13.11945, 12.66895,
    12.37225, 13.32877, 15.60949, 15.71237, 13.09488, 27.24033, 36.14561,
    18.64946, 11.44035,
  12.16347, 12.24909, 13.25913, 13.42567, 13.6665, 16.13127, 15.98522,
    13.84931, 13.76171, 14.10761, 13.5616, 12.43447, 11.71033, 14.74725,
    16.83067, 14.33796, 14.42452, 15.87991, 15.7502, 13.97995, 12.28854,
    13.20335, 16.74129, 17.91076, 15.04343, 14.57483, 23.04767, 23.43585,
    13.11815, 11.63195,
  13.92547, 14.78454, 16.44349, 17.9849, 18.46741, 16.32141, 13.2337,
    12.85859, 12.8798, 12.23959, 12.9286, 15.85478, 17.33857, 17.81616,
    17.29814, 16.81847, 17.31612, 18.06017, 17.56623, 16.28694, 15.76881,
    16.75816, 18.51625, 17.23715, 20.59716, 29.1937, 24.78269, 15.12416,
    12.35629, 10.94185,
  20.40999, 23.58187, 22.6652, 19.30426, 18.94147, 18.14126, 15.17076,
    16.52434, 17.37513, 22.75738, 26.42667, 18.5648, 16.33888, 15.88512,
    15.11566, 16.18454, 17.65777, 17.84192, 16.79675, 16.63545, 19.00948,
    19.22042, 16.61761, 14.31767, 18.87272, 24.76316, 19.2639, 12.1576,
    11.2468, 10.68618,
  32.98566, 25.88811, 25.55679, 25.65417, 24.43186, 20.67859, 24.13917,
    23.58441, 19.04994, 24.11338, 25.20544, 14.74272, 15.21601, 16.3565,
    15.45623, 16.0137, 15.71953, 15.7189, 15.33861, 15.96706, 19.13865,
    18.30417, 14.03691, 16.80045, 19.46383, 14.62683, 11.49668, 11.45257,
    11.37609, 10.86843,
  47.47915, 37.2438, 41.13511, 48.19209, 49.69049, 46.54652, 36.81486,
    21.52371, 20.63024, 20.57714, 18.04909, 12.64383, 17.25508, 19.85952,
    16.72124, 16.0948, 16.21501, 15.52145, 15.01529, 17.69905, 19.88715,
    16.58207, 13.58256, 19.33138, 21.79366, 13.41415, 11.30588, 11.63989,
    11.89354, 11.20139,
  50.0486, 65.11614, 65.28911, 68.52377, 65.03724, 55.59774, 39.65887,
    34.13476, 28.14974, 23.45511, 28.82454, 28.96516, 33.49377, 33.9533,
    29.21799, 22.10312, 16.71089, 18.18085, 19.68468, 21.30969, 19.04378,
    17.60153, 19.8623, 17.90021, 15.14351, 12.00136, 11.3811, 11.28786,
    11.73187, 11.23851,
  32.56687, 40.19466, 41.47495, 43.78913, 39.78519, 37.77114, 46.58714,
    47.2979, 37.31, 37.56648, 39.72199, 31.86736, 25.38477, 30.67225,
    33.01047, 21.01816, 19.93369, 20.06525, 21.8875, 23.74731, 21.7881,
    19.43598, 17.60438, 14.10735, 11.5017, 11.90344, 11.46334, 11.14245,
    11.18833, 10.94398,
  21.01715, 21.70517, 23.38193, 23.42876, 21.55782, 25.11123, 32.61988,
    30.08427, 27.50932, 29.59036, 28.61948, 22.14141, 17.78372, 22.65976,
    23.00323, 19.61013, 21.55742, 19.75869, 19.76864, 20.73609, 18.01358,
    15.56454, 12.78747, 12.28063, 12.2089, 11.84701, 11.49744, 11.26106,
    11.09509, 10.83165,
  19.77708, 19.64051, 19.11448, 18.00771, 17.68172, 18.98576, 20.19927,
    19.71022, 20.17861, 20.89237, 18.25068, 18.36983, 21.32574, 20.00994,
    19.78248, 20.22229, 20.384, 18.17634, 18.5867, 18.34552, 13.35411,
    13.04039, 12.69124, 12.47709, 12.15477, 11.88199, 11.43584, 11.05931,
    11.01629, 10.83312,
  17.52282, 16.97199, 15.91366, 15.89272, 16.35193, 17.33669, 18.21809,
    18.82057, 18.84667, 17.33114, 16.84135, 20.67431, 22.6266, 21.73399,
    24.17143, 22.73321, 18.92229, 16.01123, 18.09282, 17.40072, 12.79018,
    12.87781, 12.74795, 12.53106, 11.75996, 11.64609, 11.39002, 10.86981,
    10.83543, 10.74551,
  17.24469, 16.88657, 15.39577, 15.02903, 15.53936, 16.12614, 16.68597,
    16.85479, 16.13771, 15.31242, 18.139, 20.4863, 18.55854, 19.68283,
    21.35732, 20.21021, 18.8439, 17.82879, 19.56605, 18.47898, 14.80609,
    13.54888, 12.77262, 12.45566, 11.52886, 11.31513, 11.22662, 10.86115,
    10.78353, 10.70962,
  17.58907, 17.31809, 15.82932, 14.73205, 15.05552, 15.16387, 15.24496,
    15.15484, 14.77931, 16.85139, 19.52876, 17.94172, 16.27901, 16.77175,
    16.83089, 16.39488, 17.32819, 18.47985, 19.1113, 19.32807, 17.90457,
    15.39242, 12.92356, 12.50361, 11.83439, 11.31594, 11.13999, 10.89137,
    10.78003, 10.71594,
  17.05895, 17.12207, 15.86316, 14.71692, 14.68651, 14.74734, 14.61455,
    14.52551, 15.27277, 18.35895, 18.76081, 15.72135, 16.12266, 16.13884,
    15.38455, 14.76707, 14.974, 15.46399, 15.98022, 16.58555, 17.27019,
    16.66514, 14.28878, 13.08954, 12.29313, 11.60591, 11.1502, 10.89349,
    10.78277, 10.71833,
  17.64176, 16.95134, 15.7627, 15.04309, 14.85168, 14.37828, 14.48033,
    14.78573, 16.56504, 18.70885, 17.0038, 14.56779, 15.27019, 15.18209,
    14.5769, 14.11123, 13.72117, 13.62376, 14.12919, 14.23767, 15.50582,
    15.84703, 14.54966, 14.79317, 13.5794, 11.95916, 11.19733, 10.96303,
    10.79702, 10.71659,
  17.89339, 17.17156, 15.66479, 14.88036, 15.31359, 15.59091, 15.8585,
    15.76361, 17.25611, 17.84553, 15.30299, 14.09533, 14.39439, 14.27672,
    13.74632, 13.90145, 13.85899, 13.25887, 13.14367, 13.07132, 14.41125,
    14.37186, 12.91277, 14.54783, 14.80452, 12.71282, 11.39564, 11.35835,
    11.0446, 10.73915,
  17.71649, 17.1759, 16.17745, 15.9003, 16.49231, 17.01893, 18.07726,
    18.73992, 19.4195, 17.26613, 14.29774, 14.24925, 14.48451, 14.65373,
    14.31418, 14.43828, 14.67486, 13.8715, 12.97853, 13.03515, 13.471,
    13.09003, 12.39179, 12.86573, 13.93451, 14.05395, 12.71549, 11.75131,
    11.43061, 10.86959,
  17.6864, 17.6249, 16.29551, 16.2195, 17.29223, 18.06677, 18.47391,
    18.86783, 19.90801, 17.47515, 14.01099, 14.28673, 14.66431, 14.98352,
    15.00643, 15.05367, 14.7537, 14.25841, 13.48375, 13.03751, 12.95533,
    12.78205, 12.7585, 12.35383, 12.34689, 13.81782, 13.943, 12.57603,
    12.30722, 11.32929,
  17.90874, 18.82659, 18.27913, 17.79337, 17.99118, 18.19034, 18.8194,
    19.56583, 18.67001, 16.40551, 14.20955, 14.52742, 15.15517, 15.11186,
    14.6613, 14.62032, 14.20591, 13.99583, 13.77664, 13.16021, 13.12763,
    13.17275, 12.54423, 12.0135, 11.96943, 12.75788, 14.17997, 13.32818,
    12.41364, 11.3945,
  19.02847, 20.18765, 19.33341, 18.49358, 17.94163, 17.33144, 19.11411,
    19.87582, 16.92793, 14.75589, 14.56692, 15.04447, 15.34995, 14.94974,
    14.31694, 14.01056, 13.73844, 13.76526, 13.66691, 13.06816, 13.14106,
    13.98971, 13.98042, 13.40218, 13.38786, 13.61351, 15.63198, 15.2439,
    12.33247, 10.87327,
  20.10462, 20.71575, 18.57678, 18.09634, 18.23175, 17.76764, 18.79021,
    18.0055, 14.82465, 14.10802, 14.55535, 14.9501, 14.87298, 14.54107,
    14.53414, 14.21812, 13.59134, 13.44187, 13.86203, 14.26514, 14.57572,
    14.71509, 14.42148, 13.9967, 14.18723, 14.31794, 15.10065, 16.96235,
    15.02798, 11.43902,
  19.10592, 18.09368, 17.94029, 19.36025, 19.75288, 19.69773, 19.03619,
    16.16535, 14.0441, 14.20542, 13.93507, 13.67923, 13.59311, 13.71657,
    14.25369, 14.41431, 14.27586, 14.54669, 14.5582, 14.39097, 14.40917,
    13.97372, 13.13837, 12.73984, 13.1082, 13.64463, 13.79333, 14.28328,
    14.8303, 12.15781,
  18.14093, 17.74065, 18.15535, 18.70721, 18.86854, 20.02428, 19.67747,
    16.06184, 13.89389, 14.30638, 14.38083, 14.57692, 14.90724, 15.06159,
    15.19942, 15.35053, 14.78486, 14.09047, 13.74832, 13.09235, 12.61269,
    12.50781, 12.2359, 12.07467, 12.21548, 12.8319, 13.09908, 12.46401,
    12.08399, 11.1478,
  12.38614, 12.40598, 12.44023, 12.45555, 12.44252, 12.43886, 12.44037,
    12.44846, 12.46836, 12.47119, 13.12503, 13.29355, 12.51683, 12.66708,
    12.82046, 12.56911, 12.50779, 12.52254, 12.48339, 12.86185, 13.15947,
    12.80993, 12.72451, 13.05015, 13.09317, 12.65796, 14.61656, 16.40673,
    14.28728, 13.20898,
  12.6278, 12.68066, 12.52709, 12.75888, 12.63212, 12.48817, 12.50536,
    12.52492, 12.57111, 12.69663, 13.25393, 13.75198, 13.78147, 13.34375,
    13.11147, 13.12853, 12.64887, 12.6088, 12.95539, 13.5265, 13.57428,
    12.90984, 12.63668, 13.11718, 16.01287, 16.96324, 16.40595, 20.53701,
    15.84252, 14.04439,
  12.67554, 12.70743, 12.62703, 12.73707, 12.61635, 12.48734, 12.47893,
    12.54486, 12.65203, 12.75412, 12.8421, 13.26653, 13.71951, 13.94801,
    13.94121, 13.19436, 12.94562, 13.29251, 13.3458, 13.44523, 13.7069,
    14.46462, 15.1932, 14.45741, 19.0676, 23.64322, 19.11984, 20.65417,
    15.64548, 14.64385,
  12.58539, 12.5786, 12.7303, 12.80764, 12.94558, 13.32044, 13.35406,
    13.12822, 13.1242, 13.32948, 13.47458, 13.82517, 13.66422, 13.42025,
    14.20347, 14.80055, 14.39915, 13.44307, 13.156, 12.87773, 14.84519,
    16.68807, 15.73602, 19.63226, 22.74843, 21.10358, 23.04011, 19.9509,
    15.48535, 13.91428,
  12.9743, 12.65971, 12.83533, 13.07487, 13.42181, 13.72755, 13.64404,
    13.34464, 13.81652, 14.55318, 14.64014, 14.23363, 13.61062, 13.66328,
    14.50468, 15.02715, 13.80647, 12.63129, 12.68992, 16.54712, 19.26268,
    15.30894, 14.87269, 17.84293, 20.03702, 19.32267, 19.57452, 19.53793,
    19.34818, 15.03667,
  12.92141, 12.72541, 13.2927, 14.29875, 14.61601, 14.16484, 13.89493,
    13.68489, 13.6073, 13.8577, 13.63378, 14.60011, 16.2699, 16.51003,
    15.64652, 19.97026, 26.02852, 20.17412, 15.22785, 18.44601, 18.00073,
    13.92378, 14.61511, 15.51805, 18.17422, 18.38973, 18.7283, 30.43528,
    30.01297, 14.97502,
  12.75559, 12.96351, 13.83354, 15.02389, 15.44264, 14.8076, 14.7256,
    16.13047, 16.35732, 16.11173, 16.63823, 16.83388, 16.31994, 15.84776,
    19.72823, 28.0571, 27.75328, 19.20157, 16.31825, 16.57352, 15.09711,
    14.09505, 14.67156, 16.88248, 18.87835, 16.25103, 23.34778, 42.35138,
    34.39612, 13.38767,
  12.85038, 13.18985, 14.20052, 15.24007, 15.06671, 16.37031, 18.49489,
    17.40542, 16.16217, 16.34178, 16.67677, 15.73948, 14.17758, 13.89712,
    17.17142, 20.89388, 18.77802, 16.26541, 15.19961, 15.06482, 14.56647,
    14.24587, 15.32258, 17.89951, 18.10078, 15.25517, 29.38548, 41.46143,
    22.38816, 13.41069,
  13.97463, 14.10671, 15.16409, 15.39165, 15.55223, 18.45472, 18.59899,
    15.98781, 15.80824, 16.27642, 15.71697, 14.35836, 13.42552, 16.49916,
    19.19529, 16.50079, 16.33861, 18.04215, 17.93705, 16.12789, 14.15838,
    15.13496, 18.96068, 20.59378, 17.23352, 16.65376, 25.94512, 27.78685,
    15.27823, 13.61942,
  16.07635, 16.78758, 18.56469, 20.56922, 20.98908, 18.91654, 15.36172,
    14.85467, 14.88565, 14.27085, 14.71745, 17.80901, 19.44036, 20.11902,
    19.6376, 19.01299, 19.58663, 20.4811, 20.03, 18.51338, 17.89168,
    18.95901, 21.02692, 19.78041, 22.59985, 32.52539, 29.18693, 17.81686,
    14.45707, 12.82381,
  21.23481, 24.93554, 25.07797, 21.66119, 21.28575, 20.75518, 17.49446,
    18.76405, 19.81757, 24.48901, 29.13461, 21.25867, 18.6053, 18.1518,
    17.27624, 18.40782, 20.1598, 20.45053, 19.32678, 18.81007, 21.39891,
    21.80288, 19.09183, 16.35365, 21.07415, 28.34988, 23.03654, 14.24975,
    13.17376, 12.48147,
  35.94762, 28.49546, 26.85662, 26.63927, 25.74893, 21.62524, 25.89127,
    26.33713, 21.4443, 26.46812, 28.43323, 16.86574, 17.14217, 18.4727,
    17.59575, 18.35507, 18.10958, 18.11679, 17.64079, 18.19392, 21.6423,
    20.97797, 16.13148, 18.76657, 22.46376, 17.50273, 13.60995, 13.33375,
    13.25267, 12.6879,
  49.63649, 35.83937, 39.86326, 46.52135, 49.36447, 47.77706, 39.93157,
    24.35845, 23.69512, 23.32185, 20.48938, 14.19024, 19.05715, 22.17674,
    19.0671, 18.4086, 18.60391, 17.80509, 17.11975, 20.04007, 22.7001,
    18.94582, 15.51833, 21.77462, 25.71361, 15.89513, 13.18241, 13.50193,
    13.78647, 13.09214,
  52.3584, 58.45547, 58.81755, 64.33912, 65.13771, 60.10611, 44.23553,
    37.24233, 31.24945, 25.5272, 30.90544, 30.31472, 36.28701, 36.73569,
    32.3309, 24.84696, 19.08042, 20.6545, 22.33464, 24.35449, 21.97185,
    19.72237, 22.84034, 21.29601, 18.22207, 14.02782, 13.23809, 13.16844,
    13.63955, 13.16168,
  34.46657, 39.0362, 42.234, 49.35155, 51.15915, 46.07953, 49.44014,
    49.90905, 38.76044, 39.08716, 41.98013, 34.90398, 28.38306, 33.8811,
    36.67019, 23.96747, 22.61744, 22.87492, 24.9136, 26.99108, 24.51395,
    22.26882, 20.95553, 17.1131, 13.44974, 13.80736, 13.33929, 13.01866,
    13.06971, 12.82096,
  22.62264, 24.90567, 29.29271, 31.84714, 30.02246, 29.57288, 34.83381,
    31.61794, 28.53245, 31.54761, 31.13658, 24.7279, 19.73424, 25.50431,
    26.1011, 22.30817, 24.59514, 22.70514, 22.48354, 23.77912, 20.79974,
    18.47945, 15.3837, 14.45347, 14.13503, 13.76676, 13.38832, 13.13666,
    12.94862, 12.66931,
  21.00576, 21.9427, 22.3198, 20.79307, 19.05635, 19.93097, 21.50512,
    20.61466, 21.06808, 22.42597, 19.72449, 19.60279, 23.22776, 22.19451,
    22.36533, 22.95675, 23.46281, 21.05511, 21.15558, 21.66147, 16.04568,
    15.51299, 14.84196, 14.50882, 14.10918, 13.79728, 13.33577, 12.93853,
    12.85231, 12.65738,
  18.3512, 18.1354, 16.73417, 16.06135, 16.25701, 17.52277, 18.51697,
    19.11064, 19.38236, 17.89725, 17.25956, 21.75318, 24.58694, 23.64928,
    27.22182, 26.02097, 21.96959, 18.57252, 20.84707, 20.77687, 15.18524,
    15.13173, 14.7914, 14.58466, 13.72289, 13.53487, 13.29237, 12.71016,
    12.66714, 12.56377,
  17.87987, 17.39803, 15.431, 14.84305, 15.39659, 16.00545, 16.62381,
    16.93725, 16.32255, 15.24655, 18.28845, 21.59035, 19.88859, 21.56733,
    24.39994, 23.34438, 21.80014, 20.50371, 22.63407, 21.6135, 17.13373,
    15.75173, 14.83976, 14.5297, 13.47246, 13.18506, 13.11876, 12.69234,
    12.59318, 12.51521,
  18.02975, 17.41014, 15.66193, 14.3802, 14.71736, 14.89166, 15.10991,
    15.0887, 14.56532, 16.62597, 19.98143, 18.7616, 17.27275, 18.58272,
    19.34371, 19.08353, 20.17594, 21.55453, 22.16369, 22.27967, 20.45781,
    17.86914, 15.05528, 14.55143, 13.78106, 13.20625, 13.00919, 12.73005,
    12.58871, 12.51616,
  17.20776, 16.99868, 15.60988, 14.33819, 14.35652, 14.52714, 14.45469,
    14.24516, 14.89449, 18.32325, 19.38292, 16.27272, 17.25559, 18.00631,
    17.67671, 17.26222, 17.66424, 18.2547, 18.59056, 19.27425, 19.99671,
    19.41059, 16.52791, 15.18378, 14.26433, 13.52526, 13.01771, 12.73268,
    12.59303, 12.52104,
  17.77033, 16.7494, 15.5133, 14.74138, 14.65112, 14.15579, 14.16401,
    14.34817, 16.29754, 18.94338, 17.49263, 15.10358, 16.54367, 17.08295,
    16.84025, 16.5465, 16.20375, 15.97115, 16.47273, 16.65643, 18.00913,
    18.65364, 16.75777, 17.05156, 15.7298, 13.96402, 13.06773, 12.8004,
    12.60227, 12.52103,
  18.02516, 17.01193, 15.4726, 14.64627, 15.15289, 15.33599, 15.51654,
    15.41215, 17.21021, 18.25478, 15.68581, 14.75981, 15.69975, 16.13777,
    15.94158, 16.23699, 16.20245, 15.50955, 15.37572, 15.27298, 16.74346,
    17.03591, 14.98581, 16.83056, 17.13993, 14.83265, 13.25663, 13.22711,
    12.87826, 12.54475,
  17.87447, 17.09663, 16.09415, 15.7378, 16.31161, 16.74704, 17.9926,
    18.95192, 19.93718, 17.84549, 14.64481, 14.99241, 15.7984, 16.5162,
    16.48475, 16.71778, 17.04231, 16.21674, 15.16217, 15.14157, 15.77258,
    15.41935, 14.41549, 15.03527, 16.17869, 16.2142, 14.72722, 13.66615,
    13.30155, 12.6974,
  17.80796, 17.65619, 16.20029, 15.96256, 17.10739, 18.08519, 18.7651,
    19.45483, 20.70279, 18.25504, 14.43749, 15.12008, 15.99515, 16.84552,
    17.17938, 17.44747, 17.2206, 16.64255, 15.6796, 15.15132, 15.11401,
    14.87177, 14.83751, 14.46373, 14.38178, 15.89041, 16.09177, 14.57654,
    14.21358, 13.2607,
  18.07526, 18.88542, 18.21193, 17.66713, 17.9988, 18.53409, 19.45255,
    20.46157, 19.51501, 17.18977, 14.68349, 15.34681, 16.46603, 16.95252,
    16.84478, 17.05593, 16.63333, 16.27107, 15.98512, 15.25386, 15.2107,
    15.30358, 14.64875, 13.99602, 13.8786, 14.73089, 16.25583, 15.46237,
    14.35635, 13.36226,
  19.22499, 20.15455, 19.35159, 18.51672, 18.14189, 17.74944, 20.00789,
    21.17354, 17.81449, 15.26224, 15.01014, 15.83606, 16.71323, 16.81955,
    16.50568, 16.33903, 16.02779, 15.97317, 15.86772, 15.15303, 15.21439,
    16.12845, 16.13442, 15.41204, 15.35863, 15.65514, 17.75614, 17.54186,
    14.3455, 12.74502,
  20.46353, 21.06059, 18.57303, 18.22897, 18.63804, 18.35018, 19.7804,
    19.22523, 15.4223, 14.38437, 14.95687, 15.75852, 16.25553, 16.4114,
    16.7262, 16.52012, 15.81505, 15.60399, 15.9767, 16.35276, 16.74218,
    17.01014, 16.68237, 16.15759, 16.27388, 16.50472, 17.36796, 19.30124,
    17.34853, 13.39212,
  19.42471, 18.2562, 18.08637, 20.09799, 20.69392, 20.63854, 20.16209,
    17.03131, 14.30944, 14.4318, 14.32346, 14.42347, 14.84249, 15.43908,
    16.36824, 16.68951, 16.49494, 16.74993, 16.77011, 16.56518, 16.65222,
    16.21736, 15.26988, 14.80382, 15.18458, 15.78739, 16.00784, 16.56751,
    17.09225, 14.27837,
  18.59268, 18.13115, 18.89378, 19.90512, 20.14197, 21.29611, 20.88043,
    16.78796, 14.1214, 14.62931, 14.84358, 15.33879, 16.1384, 16.80369,
    17.29564, 17.60443, 17.06985, 16.31541, 15.91473, 15.17522, 14.63926,
    14.5119, 14.20843, 14.0246, 14.21467, 14.87766, 15.2205, 14.57008,
    14.10359, 13.07768,
  16.02967, 16.06887, 16.08885, 16.1124, 16.09992, 16.09474, 16.09261,
    16.1099, 16.14351, 16.16809, 16.94901, 17.20984, 16.20892, 16.37791,
    16.58067, 16.25297, 16.16627, 16.18898, 16.15485, 16.61655, 17.01634,
    16.59227, 16.52033, 16.90163, 16.93875, 16.47986, 18.67155, 21.1173,
    18.50814, 17.21791,
  16.30076, 16.41878, 16.19153, 16.47288, 16.32584, 16.13902, 16.16682,
    16.19341, 16.25613, 16.44159, 17.05581, 17.64204, 17.73751, 17.21362,
    16.86443, 16.92857, 16.32377, 16.29345, 16.73095, 17.42069, 17.45334,
    16.66218, 16.34604, 17.00444, 20.39675, 22.2352, 21.16407, 26.53119,
    20.41142, 18.24201,
  16.3688, 16.40202, 16.30965, 16.42279, 16.28075, 16.14327, 16.13086,
    16.21308, 16.35268, 16.47672, 16.60712, 17.10195, 17.59051, 17.88433,
    17.93113, 17.00147, 16.70974, 17.17801, 17.22185, 17.32885, 17.68047,
    18.69984, 19.60312, 18.97127, 24.04523, 30.22537, 24.91275, 26.87949,
    20.21615, 19.02218,
  16.28577, 16.25737, 16.41285, 16.5467, 16.71158, 17.17203, 17.23244,
    16.94197, 16.9208, 17.15963, 17.34997, 17.77221, 17.64149, 17.26505,
    18.22754, 19.01908, 18.60979, 17.38418, 16.95938, 16.71865, 19.13536,
    21.48546, 20.30729, 24.86822, 28.70938, 26.66435, 30.15957, 25.86121,
    20.09577, 18.07584,
  16.76082, 16.34295, 16.55228, 16.84276, 17.27169, 17.61776, 17.51307,
    17.196, 17.75638, 18.77369, 18.99625, 18.33449, 17.4634, 17.70689,
    18.72375, 19.18618, 17.86159, 16.36259, 16.50879, 21.10966, 24.65023,
    19.6883, 19.27859, 22.48066, 25.01494, 24.49234, 25.01426, 25.73733,
    25.56409, 19.46597,
  16.64204, 16.43047, 17.14067, 18.36448, 18.82664, 18.29823, 17.84589,
    17.62007, 17.47788, 17.78157, 17.60624, 18.75484, 20.93559, 21.1476,
    20.47806, 25.06319, 32.13528, 25.70155, 19.87465, 23.42852, 22.8162,
    17.95024, 18.77693, 19.98586, 22.89569, 23.34512, 23.4024, 37.22515,
    37.94833, 19.36456,
  16.47211, 16.74883, 17.80364, 19.20468, 19.84172, 19.17481, 18.84721,
    20.68367, 21.03134, 20.73962, 21.41667, 21.68145, 20.91396, 20.46006,
    24.79178, 33.9114, 33.51577, 24.17661, 20.94209, 21.21853, 19.35761,
    18.07673, 18.80478, 21.46252, 23.78771, 21.10581, 27.8788, 48.55298,
    42.04206, 17.56467,
  16.57651, 17.02459, 18.24028, 19.51906, 19.35457, 20.88434, 23.57996,
    22.27544, 20.61708, 20.91987, 21.28845, 20.22757, 18.27851, 18.15942,
    21.93492, 26.03993, 23.48561, 20.98321, 19.47563, 19.25229, 18.60798,
    18.20948, 19.58237, 22.67168, 22.9339, 20.09191, 34.75392, 49.20396,
    27.60403, 17.45368,
  18.0535, 18.28666, 19.4169, 19.64362, 19.92857, 23.75793, 24.00068,
    20.40591, 20.35323, 20.92337, 20.22509, 18.5019, 17.45306, 21.15066,
    24.8459, 21.56173, 20.84135, 22.90457, 22.83336, 20.62159, 18.10893,
    19.41752, 24.0492, 26.1135, 21.83669, 21.5867, 31.67568, 34.55009,
    19.83373, 17.56283,
  20.31203, 20.80294, 23.3757, 26.81669, 26.8324, 24.16486, 19.67479,
    18.97207, 18.97214, 18.38789, 18.8538, 22.64268, 24.65762, 25.4626,
    24.6631, 23.9069, 24.74595, 25.81631, 25.12971, 23.11821, 22.56011,
    23.85147, 26.18474, 24.91196, 28.24317, 40.16442, 36.85014, 22.73609,
    18.44351, 16.58051,
  27.80922, 34.51656, 34.74273, 27.33135, 27.12307, 26.4189, 23.18865,
    24.4037, 25.78541, 29.6845, 35.45863, 26.74344, 23.78418, 23.18929,
    22.16026, 23.56196, 25.78965, 26.12572, 24.62013, 23.39408, 26.37127,
    26.92761, 23.78938, 20.72921, 26.04531, 34.13572, 28.35281, 18.15496,
    17.00322, 16.1409,
  46.19397, 37.93438, 34.11341, 31.00625, 31.35215, 26.04201, 30.73492,
    31.39291, 26.85969, 32.25204, 33.93442, 21.35942, 21.8663, 23.41387,
    22.49095, 23.59149, 23.34988, 23.34652, 22.56051, 22.92193, 26.84916,
    25.99863, 20.35858, 23.1633, 28.02806, 22.52579, 17.61177, 17.12132,
    17.04984, 16.3926,
  60.49564, 46.10694, 48.33363, 54.49154, 56.69999, 53.83931, 47.77995,
    40.54891, 46.60221, 33.90912, 24.38049, 19.02265, 24.73986, 27.48509,
    24.96289, 23.39241, 23.77768, 22.78338, 21.70348, 25.04336, 28.30903,
    23.5271, 19.75525, 26.39957, 31.48491, 20.20223, 16.94027, 17.34189,
    17.65108, 16.90118,
  67.91483, 58.64676, 60.93524, 67.08909, 70.33176, 69.88632, 61.05404,
    59.07532, 49.46902, 33.40963, 37.13403, 39.11411, 44.84207, 45.8269,
    40.36209, 30.29892, 24.38262, 26.33459, 28.60002, 31.16598, 28.01331,
    24.22245, 28.36321, 26.47511, 22.8125, 18.01079, 17.02865, 16.96018,
    17.46603, 16.98716,
  49.82723, 61.7519, 73.15276, 78.93022, 78.7473, 69.1861, 66.53465, 68.267,
    48.1172, 47.19341, 52.60682, 43.86676, 36.27337, 42.70788, 44.42813,
    30.55014, 28.91178, 29.48763, 32.11523, 34.19918, 29.7848, 27.32014,
    26.18347, 21.81201, 17.40089, 17.69589, 17.14927, 16.79751, 16.82536,
    16.56824,
  36.77637, 47.35484, 55.95423, 55.55074, 48.04388, 46.19539, 49.98164,
    39.73696, 36.87487, 41.23067, 41.38468, 32.84452, 26.1944, 32.53898,
    32.44315, 28.68799, 31.47782, 29.25873, 28.31488, 29.64694, 25.50427,
    22.9996, 19.91164, 18.63805, 18.07024, 17.64608, 17.20206, 16.94095,
    16.7047, 16.37923,
  29.25567, 30.55166, 31.062, 28.14672, 25.15372, 28.12963, 30.46373,
    26.47173, 28.72075, 30.44887, 26.12525, 25.27119, 29.05356, 27.50318,
    28.21576, 29.0241, 30.10553, 26.99717, 26.49771, 27.93545, 20.6324,
    19.80338, 18.97067, 18.62063, 18.08242, 17.67955, 17.17614, 16.71467,
    16.58864, 16.36851,
  23.01245, 22.87465, 20.81631, 19.69523, 20.26088, 22.15337, 23.22135,
    24.01328, 24.37567, 22.37295, 21.14939, 26.42733, 30.05909, 28.57442,
    34.12621, 32.95176, 28.05672, 23.54613, 26.26867, 26.7312, 19.4204,
    19.47149, 18.9594, 18.71285, 17.63692, 17.38855, 17.15066, 16.45303,
    16.37704, 16.26083,
  21.98815, 21.37475, 18.7328, 17.89792, 18.59658, 19.29906, 20.11931,
    20.44691, 19.58732, 18.15383, 21.6088, 25.71784, 23.72462, 26.00263,
    30.66778, 29.38248, 27.57678, 25.74914, 28.61616, 27.46952, 21.82011,
    20.27531, 19.13141, 18.69312, 17.34962, 17.00769, 16.93794, 16.42294,
    16.30054, 16.19845,
  21.68257, 20.73141, 18.52073, 16.91972, 17.37805, 17.62652, 17.86559,
    17.83261, 17.16738, 19.48985, 23.55025, 21.96476, 20.19209, 22.33419,
    23.93585, 24.1407, 25.70741, 27.53686, 28.19844, 28.31309, 25.78789,
    22.79216, 19.45836, 18.73252, 17.71346, 17.03841, 16.80307, 16.47079,
    16.28226, 16.19991,
  20.34079, 19.97411, 18.2092, 16.63335, 16.69052, 16.90778, 16.82928,
    16.5651, 17.31506, 21.33492, 22.68967, 18.75074, 20.07445, 21.38266,
    21.50088, 21.65717, 22.65172, 23.75686, 24.06638, 24.85613, 25.70036,
    25.20125, 21.16711, 19.48273, 18.23906, 17.41865, 16.81449, 16.48027,
    16.28795, 16.20592,
  21.07701, 19.46643, 17.97333, 16.98443, 16.9402, 16.33505, 16.36352,
    16.5371, 18.87964, 22.11286, 20.34352, 17.28576, 19.26781, 20.3012,
    20.52385, 20.71776, 20.79172, 20.74347, 21.4234, 21.79924, 23.40324,
    24.33805, 21.41549, 21.74586, 20.11114, 18.02636, 16.89956, 16.57834,
    16.30123, 16.20753,
  21.3324, 19.67886, 17.85905, 16.78777, 17.48953, 17.70411, 17.84614,
    17.64879, 19.85358, 21.30703, 18.06282, 16.91247, 18.2845, 19.21844,
    19.52246, 20.39173, 20.75289, 20.08534, 20.01409, 20.01928, 21.58069,
    22.08697, 19.43173, 21.65768, 21.95338, 19.12419, 17.08698, 17.06646,
    16.63564, 16.24114,
  21.17007, 19.69984, 18.60155, 18.16524, 18.88761, 19.24858, 20.82521,
    22.32311, 23.55139, 20.82827, 16.8515, 17.3425, 18.50515, 19.72758,
    20.21358, 20.98805, 21.74678, 20.94458, 19.72371, 19.82955, 20.69802,
    20.12271, 18.65696, 19.61831, 20.91946, 20.75861, 18.95233, 17.597,
    17.10749, 16.435,
  20.80739, 20.72717, 18.78729, 18.26616, 19.74682, 21.1641, 22.11503,
    23.1388, 24.3765, 21.44313, 16.72036, 17.66117, 18.83745, 20.20535,
    21.06538, 21.95994, 22.07537, 21.50901, 20.31513, 19.64509, 19.71869,
    19.29107, 19.23564, 18.94584, 18.62934, 20.2756, 20.4681, 18.63213,
    18.12164, 17.13864,
  21.23393, 22.50327, 21.44799, 20.61755, 21.05853, 21.9129, 23.19913,
    24.56684, 23.04386, 20.39927, 17.21707, 18.05088, 19.45164, 20.39642,
    20.74324, 21.57078, 21.47853, 21.0627, 20.58503, 19.53728, 19.52042,
    19.75552, 19.06273, 18.13904, 17.81922, 18.84706, 20.48987, 19.7037,
    18.32551, 17.28753,
  22.58593, 23.85676, 22.8685, 21.44888, 21.23815, 21.11901, 24.20642,
    25.74449, 21.22231, 18.18566, 17.75247, 18.70858, 19.79521, 20.22264,
    20.36027, 20.73509, 20.68684, 20.65037, 20.4078, 19.35592, 19.55834,
    20.71131, 20.65644, 19.59202, 19.43556, 19.86297, 22.15565, 22.11762,
    18.36371, 16.50672,
  24.71173, 26.55549, 21.56039, 20.82556, 21.7229, 21.77393, 23.72918,
    23.3385, 18.47593, 17.14408, 17.79008, 18.71243, 19.32977, 19.73025,
    20.60635, 20.93702, 20.35443, 20.1497, 20.41965, 20.64486, 21.33498,
    21.92895, 21.44003, 20.61923, 20.53212, 20.93777, 21.97595, 24.02732,
    21.85562, 17.28603,
  23.29004, 21.88396, 21.02653, 24.95791, 25.33624, 24.29848, 24.22169,
    20.59412, 17.11307, 17.22549, 17.10847, 17.11711, 17.59456, 18.52172,
    20.12119, 21.06108, 21.09591, 21.45748, 21.38904, 21.02471, 21.29913,
    20.89991, 19.69801, 19.02024, 19.40207, 20.15555, 20.49538, 21.16945,
    21.59366, 18.4281,
  21.95408, 21.08171, 22.97301, 25.911, 25.52043, 25.75599, 25.26169,
    20.3681, 16.90278, 17.54031, 17.7085, 18.13255, 19.02187, 20.03096,
    21.12427, 22.04691, 21.79717, 21.02665, 20.43407, 19.45463, 18.85042,
    18.61683, 18.23595, 18.01189, 18.29341, 19.06653, 19.49364, 18.80084,
    18.19018, 16.97288,
  19.05124, 19.1225, 19.20192, 19.24692, 19.21365, 19.22092, 19.22475,
    19.26466, 19.34313, 19.59927, 21.04419, 21.59453, 19.54951, 19.8916,
    20.24572, 19.55058, 19.36028, 19.44521, 19.48559, 20.16174, 20.83842,
    20.38664, 20.68591, 21.50844, 22.20997, 22.64849, 26.64117, 30.78457,
    24.0382, 21.14089,
  19.67909, 19.93531, 19.45145, 19.95244, 19.65491, 19.31247, 19.41407,
    19.51769, 19.71405, 20.16757, 21.10077, 22.11393, 22.55911, 21.56516,
    20.67393, 20.91644, 19.78176, 19.91825, 20.82882, 21.89604, 21.7486,
    20.73821, 20.97984, 23.84459, 30.81136, 35.22363, 31.79956, 38.8187,
    26.66709, 22.66761,
  19.67136, 19.71602, 19.5837, 19.69507, 19.45562, 19.32661, 19.39288,
    19.57887, 19.82611, 20.0204, 20.31359, 21.16857, 21.92703, 22.58416,
    22.80214, 21.06063, 20.78295, 21.66781, 21.60414, 22.01479, 23.6467,
    27.0247, 29.52073, 30.49967, 39.26069, 47.88944, 39.56177, 39.13107,
    26.53873, 24.11637,
  19.57398, 19.58852, 19.86723, 20.17797, 20.57389, 21.42621, 21.5182,
    21.0039, 21.04395, 21.65338, 22.20516, 22.64494, 22.36939, 21.69804,
    23.62511, 25.26966, 24.3137, 21.85826, 21.75846, 23.13753, 29.03565,
    33.89991, 31.68587, 38.97559, 46.81794, 41.83936, 47.424, 36.68439,
    26.35176, 22.2805,
  20.47296, 19.74567, 20.37786, 21.07658, 21.79829, 22.06583, 21.8506,
    21.69059, 22.95586, 24.46378, 24.03975, 22.95001, 22.14129, 22.87791,
    24.23649, 24.52555, 23.15677, 21.85798, 23.73615, 31.93714, 37.54854,
    29.60195, 29.99117, 34.0316, 36.20448, 35.97651, 35.57224, 38.99561,
    36.3938, 23.59328,
  20.23635, 20.55261, 22.36991, 24.71371, 24.67844, 23.06437, 22.76069,
    22.22183, 21.91728, 22.10869, 22.3263, 25.28063, 30.13851, 30.86833,
    33.64924, 40.2486, 46.07467, 39.52854, 31.53616, 35.55318, 33.09423,
    25.93267, 27.92615, 30.51102, 33.26246, 33.87638, 38.16297, 58.4621,
    53.46685, 24.69302,
  20.52841, 21.7447, 23.95484, 26.21729, 25.92403, 24.33323, 25.96947,
    30.30368, 31.21384, 30.95558, 32.05798, 31.49735, 29.67468, 30.73806,
    38.05302, 48.7914, 45.43074, 36.20504, 31.13617, 30.99804, 27.65208,
    25.60645, 27.63505, 33.03418, 37.55693, 38.50403, 49.62148, 64.92347,
    54.92495, 21.55736,
  20.86614, 22.3867, 24.90319, 27.03364, 26.42424, 29.35196, 35.58061,
    33.64683, 29.9453, 30.76361, 30.18469, 27.66281, 25.234, 27.24512,
    32.31457, 36.16472, 33.41048, 31.6556, 27.25036, 26.81427, 25.46496,
    25.24256, 28.79368, 34.63302, 36.2477, 36.68254, 51.78837, 62.51634,
    37.93975, 21.32659,
  23.47805, 24.24039, 26.34885, 27.27831, 29.25773, 34.56627, 32.6115,
    28.87878, 29.3496, 29.07756, 27.27476, 24.6545, 24.79871, 33.03135,
    40.15206, 32.53639, 30.42634, 33.92693, 33.77414, 29.4821, 25.05442,
    28.89744, 37.82013, 41.4288, 33.98431, 36.50015, 49.4302, 49.01004,
    27.24757, 21.43614,
  27.94145, 32.81084, 35.41281, 38.24659, 39.37524, 35.95871, 24.791,
    24.53847, 23.76543, 23.9825, 27.41773, 36.36079, 40.28699, 40.04024,
    37.05708, 35.7967, 37.83066, 39.38792, 35.35296, 31.05468, 31.6136,
    33.87958, 36.8969, 37.92456, 47.24928, 61.34198, 53.67296, 30.18263,
    22.18972, 19.69001,
  43.45681, 48.60802, 49.86346, 47.2379, 46.5757, 37.40036, 30.78452,
    34.22825, 38.71846, 45.70075, 53.87766, 39.08203, 33.52802, 32.50773,
    31.79486, 34.05587, 37.02415, 36.47581, 33.17984, 31.21397, 34.84663,
    35.84544, 31.47393, 29.33143, 36.60155, 43.07398, 33.83146, 21.10379,
    20.27357, 19.13877,
  64.59042, 51.08192, 51.68837, 52.58637, 50.10998, 39.64452, 47.81746,
    49.56938, 44.97322, 46.96141, 43.63674, 29.21906, 30.79171, 33.24357,
    32.75818, 34.30347, 33.50199, 32.41045, 30.97603, 32.25329, 35.65738,
    33.42638, 26.63826, 31.39487, 37.2036, 27.92876, 20.85527, 20.48023,
    20.42563, 19.52657,
  79.48306, 67.62137, 80.13838, 87.97651, 88.40005, 81.3375, 67.69054,
    49.69926, 51.29456, 40.99577, 32.87802, 28.48271, 36.45485, 41.70903,
    38.78957, 34.76431, 34.05664, 31.9366, 30.53903, 37.56459, 40.41918,
    29.75823, 26.97649, 34.18341, 38.42797, 23.93112, 20.10646, 20.92089,
    21.24084, 20.23029,
  89.08198, 104.166, 104.4577, 105.1663, 96.5012, 87.79488, 78.18094,
    71.42153, 57.01564, 47.43935, 58.57513, 59.43409, 65.94758, 67.05823,
    59.24969, 44.49146, 35.46514, 38.06579, 41.66488, 44.3622, 38.56314,
    32.16805, 37.06438, 32.00084, 25.96601, 21.53363, 20.47557, 20.3292,
    20.87837, 20.28639,
  84.13741, 83.68442, 86.17582, 82.14304, 71.62376, 70.74361, 83.69592,
    80.89436, 69.37976, 73.41747, 76.24453, 65.69887, 59.4071, 65.00423,
    62.74451, 46.24937, 44.43074, 46.97386, 51.65842, 51.75757, 41.77658,
    39.09556, 34.10193, 25.08594, 20.83022, 21.28317, 20.57821, 20.07883,
    20.04363, 19.69701,
  75.69566, 73.7872, 71.38893, 64.13729, 60.7124, 66.39319, 82.52753,
    83.71163, 62.35131, 64.89626, 62.44555, 52.16439, 46.30555, 53.39343,
    50.24501, 46.75838, 49.45932, 46.53662, 46.38877, 46.82902, 34.49232,
    29.58675, 25.16387, 22.43402, 21.85341, 21.2268, 20.55745, 20.21529,
    19.86308, 19.4641,
  61.61988, 57.84704, 51.68173, 50.64565, 50.38138, 50.70803, 59.00863,
    64.3726, 49.62062, 50.59569, 45.2093, 43.01833, 49.0724, 47.83164,
    47.08752, 47.39418, 46.92282, 41.96461, 42.42517, 41.86788, 26.07204,
    23.40129, 22.91898, 23.11511, 21.9771, 21.24513, 20.53967, 19.86798,
    19.68323, 19.45277,
  45.6623, 41.95108, 37.49377, 38.72341, 40.90252, 44.81438, 48.0475,
    47.28427, 42.44717, 39.00779, 39.47085, 48.1243, 52.17236, 52.0618,
    56.65889, 51.56105, 42.47788, 36.77102, 41.10334, 37.61752, 23.62319,
    24.44592, 24.14008, 23.4582, 21.16672, 20.79826, 20.51791, 19.51524,
    19.41367, 19.28796,
  39.02457, 37.14729, 33.11084, 32.2551, 36.6375, 39.95913, 38.63168,
    35.98701, 33.37833, 32.37603, 39.53678, 47.45175, 44.68855, 48.67294,
    50.49334, 43.18559, 40.73487, 42.2226, 45.22553, 39.75401, 29.0539,
    27.39723, 25.17319, 23.26298, 20.67733, 20.32872, 20.18413, 19.48037,
    19.31913, 19.21274,
  36.21835, 36.35328, 32.25102, 29.84521, 33.25014, 33.58401, 30.77475,
    28.91789, 28.46523, 35.25988, 44.3021, 41.56807, 39.80725, 41.71079,
    39.43406, 35.21259, 36.73777, 42.10732, 44.18929, 43.43971, 38.01471,
    31.48256, 25.57645, 23.24679, 21.27032, 20.43277, 20.04256, 19.5738,
    19.3136, 19.22774,
  34.73002, 35.21677, 30.37176, 28.06996, 29.40828, 28.80599, 26.72001,
    26.3896, 29.10425, 38.2617, 42.53119, 35.62246, 37.71088, 36.21384,
    33.2243, 31.73798, 33.44876, 37.28386, 39.28774, 39.73333, 37.27728,
    33.82095, 28.05223, 24.35166, 21.91771, 20.97055, 20.07829, 19.62206,
    19.34296, 19.24027,
  35.48989, 33.70529, 29.58791, 27.7788, 27.64949, 25.439, 25.44114,
    26.89728, 32.77069, 39.79511, 37.08188, 31.75711, 33.61264, 31.39267,
    29.50467, 29.69417, 31.30573, 33.80679, 35.05111, 33.76089, 32.82804,
    32.324, 29.38801, 28.53446, 25.41053, 22.11539, 20.24824, 19.7919,
    19.36982, 19.24632,
  34.67907, 33.21796, 28.18857, 26.12556, 27.37652, 27.76898, 28.62806,
    29.49961, 34.93821, 38.15302, 31.2739, 28.47985, 28.89743, 27.87126,
    27.24413, 29.15298, 31.87017, 32.00058, 31.12107, 29.63642, 29.76497,
    29.47989, 27.20837, 29.22053, 28.77995, 23.99464, 20.5964, 20.5777,
    19.85483, 19.29787,
  34.42517, 31.97507, 29.40521, 29.0336, 30.63802, 31.37659, 33.98345,
    35.16171, 38.81102, 36.37277, 27.6939, 27.23089, 27.84247, 28.37957,
    28.86554, 31.28749, 33.96754, 32.63934, 29.64249, 28.50331, 27.94918,
    26.9992, 26.19012, 27.18266, 28.07997, 26.85237, 23.67893, 21.34089,
    20.48027, 19.59514,
  32.46647, 33.97903, 28.99861, 28.58622, 31.57215, 33.32518, 34.72353,
    35.95783, 40.0924, 36.07031, 26.06882, 27.07509, 28.52721, 30.19876,
    31.78572, 34.26458, 34.49109, 32.59125, 29.11201, 26.25756, 26.45537,
    26.98265, 26.44905, 25.02692, 23.97869, 25.6109, 25.52571, 22.78171,
    21.88721, 20.62701,
  34.15518, 37.36125, 33.77031, 32.46021, 33.46346, 33.91385, 35.45315,
    38.32178, 39.39779, 32.92688, 26.45822, 28.11638, 30.76953, 32.46415,
    33.02309, 34.1545, 33.00746, 30.85393, 27.92714, 24.91813, 26.62456,
    28.01205, 25.30506, 22.52746, 21.77208, 23.32248, 25.3637, 24.3174,
    22.16077, 20.82917,
  37.70788, 40.9133, 37.604, 34.54713, 34.69298, 33.72752, 36.63579,
    38.56111, 35.13404, 28.74611, 27.75391, 30.4312, 32.91888, 33.50869,
    32.96515, 32.32184, 30.78898, 29.13421, 26.79453, 24.50603, 26.58343,
    28.99024, 27.36866, 24.6343, 23.95306, 24.90075, 27.77809, 27.63666,
    22.28058, 19.70939,
  41.51402, 43.90284, 36.38585, 34.39807, 36.95596, 36.70089, 38.43205,
    37.01393, 29.44671, 27.43201, 29.37315, 32.19617, 33.73678, 33.38417,
    32.98248, 31.60418, 29.15715, 27.61542, 26.49403, 26.39676, 29.46032,
    31.25743, 28.57526, 26.22537, 25.48613, 26.44633, 27.80782, 30.18687,
    27.16506, 20.84329,
  36.88869, 32.63787, 32.8387, 37.81121, 40.40841, 42.4249, 40.53943,
    33.06459, 26.81311, 28.29065, 29.55019, 30.48836, 31.06794, 31.1991,
    31.62087, 31.0043, 29.98758, 29.81894, 28.25922, 27.04316, 28.72897,
    28.20429, 25.31488, 23.77264, 24.11757, 25.32377, 25.91223, 26.59104,
    26.61366, 22.49707,
  33.00249, 31.86545, 35.76114, 38.22722, 38.01127, 41.19351, 42.06051,
    32.23661, 26.60302, 29.56712, 31.42127, 32.75894, 33.29762, 33.2058,
    33.08093, 32.97601, 31.31042, 28.9162, 26.73549, 24.70311, 24.06078,
    23.2369, 22.42531, 22.09048, 22.60835, 23.66438, 24.21295, 23.31924,
    22.13557, 20.32306,
  23.04235, 23.40174, 23.80371, 24.21863, 24.37602, 24.7102, 25.13758,
    25.71623, 26.52249, 27.92029, 30.52043, 30.71325, 26.14113, 27.15641,
    27.56828, 26.43181, 26.90651, 28.42725, 30.44519, 33.68394, 35.80411,
    34.73718, 36.29309, 39.88053, 43.19749, 44.67674, 51.06707, 54.25936,
    33.29221, 26.72062,
  25.06629, 25.78339, 24.84538, 26.23255, 25.67416, 25.45317, 26.20373,
    26.88271, 27.851, 29.12923, 31.04438, 33.49434, 34.66614, 31.86915,
    30.33617, 32.04289, 31.26402, 34.16947, 37.97169, 41.35917, 42.4498,
    43.28716, 46.40234, 54.15329, 61.97411, 58.73767, 52.56293, 56.48828,
    35.02244, 28.76695,
  22.70165, 22.92537, 23.27619, 23.743, 24.03985, 24.55621, 25.07998,
    25.86077, 26.87974, 28.04753, 29.59932, 32.23238, 35.08126, 38.50951,
    41.07419, 39.82354, 42.98216, 47.64794, 51.18118, 57.02905, 65.44537,
    73.7661, 76.77282, 77.26734, 78.0036, 72.39857, 65.89027, 54.24887,
    35.45094, 30.96976,
  24.47873, 25.39007, 27.27125, 29.36888, 31.25763, 33.44305, 33.77588,
    33.37481, 34.58142, 36.46751, 37.81607, 39.62699, 41.48634, 43.57812,
    51.27555, 56.60042, 55.39534, 54.08859, 60.44518, 67.78761, 78.35522,
    81.71105, 76.19505, 82.49866, 82.29161, 79.19621, 71.84145, 52.59431,
    35.40805, 27.65056,
  29.15494, 28.55131, 31.21607, 33.00011, 34.41993, 34.22833, 34.07224,
    34.9789, 37.99023, 40.48538, 40.21973, 42.25167, 45.23501, 49.99605,
    55.08242, 59.00677, 58.84904, 56.44473, 61.98653, 71.73297, 74.47664,
    63.48108, 65.19327, 73.325, 79.68336, 78.75978, 71.20723, 75.39453,
    64.06377, 35.92482,
  30.13079, 32.77755, 36.73376, 40.92215, 40.20228, 38.2314, 40.42065,
    42.80351, 45.39999, 51.06014, 59.24466, 72.21736, 85.47101, 85.28086,
    88.73049, 93.63085, 93.84032, 84.75101, 72.65337, 72.63036, 64.67899,
    57.3015, 64.21672, 71.82355, 79.68449, 79.63638, 76.5827, 89.71296,
    75.28654, 33.85107,
  34.73627, 40.11494, 46.3798, 53.3013, 57.42851, 62.55012, 72.84062,
    83.38084, 86.21492, 86.03892, 85.98578, 79.8422, 70.25082, 71.05862,
    73.30144, 75.58235, 75.44401, 68.92664, 59.8937, 61.18016, 58.30666,
    58.71931, 64.93454, 73.69353, 75.97446, 67.7247, 70.46741, 79.88215,
    63.21742, 26.02238,
  43.17111, 51.10923, 59.24606, 67.31609, 71.08995, 79.93612, 85.76527,
    70.20662, 59.63948, 58.99321, 54.17742, 48.82677, 44.73042, 46.58796,
    50.24129, 55.97257, 59.70908, 59.50706, 53.22299, 54.61052, 54.73073,
    58.20006, 66.50078, 72.60186, 68.29939, 64.1457, 74.70975, 74.40479,
    49.67276, 26.97828,
  56.57089, 61.01908, 65.77586, 67.77838, 66.86383, 69.09012, 59.16923,
    53.10426, 54.7921, 54.85664, 53.80665, 53.51299, 57.92889, 72.05318,
    81.32964, 67.07269, 69.7364, 77.19788, 76.33398, 68.16542, 65.37605,
    78.54646, 92.1172, 91.20103, 76.66092, 82.87823, 82.72042, 66.25396,
    35.27206, 26.69651,
  79.80809, 86.90959, 82.98681, 85.91285, 77.75557, 65.99884, 48.81997,
    57.57419, 61.27782, 71.82971, 83.59995, 95.68359, 94.92961, 91.28217,
    85.4893, 93.10012, 99.04186, 97.5459, 90.96001, 87.72776, 95.26477,
    94.09241, 89.59888, 79.79132, 85.68065, 96.23021, 77.69066, 43.49186,
    26.59852, 23.24878,
  103.0791, 96.43726, 95.80543, 85.97677, 96.6688, 97.90347, 95.61059,
    102.0378, 108.6556, 111.2016, 100.8765, 74.65411, 71.76147, 73.25197,
    77.08319, 84.00294, 88.93371, 87.86418, 84.25249, 83.64436, 93.58475,
    88.27136, 67.47094, 59.65962, 65.7357, 63.60204, 42.7945, 26.71789,
    25.32861, 22.94992,
  108.4765, 93.04886, 104.6464, 112.7408, 110.4284, 95.23538, 97.79871,
    91.22177, 81.02064, 69.51907, 62.09752, 58.0952, 65.49175, 72.3774,
    75.30979, 76.01086, 74.11366, 72.47574, 69.25561, 70.53147, 78.79487,
    71.63137, 54.04399, 62.65248, 64.95787, 44.64017, 25.92381, 28.03912,
    26.36446, 24.13678,
  121.6516, 122.4647, 125.6852, 126.4564, 124.8161, 120.0054, 95.43832,
    83.6984, 85.94566, 65.56248, 64.66959, 67.41205, 79.22517, 87.89882,
    83.76665, 71.01154, 71.63686, 68.07865, 65.63898, 71.74374, 74.6382,
    63.1772, 55.55556, 54.99037, 51.20921, 36.33221, 27.67516, 29.64414,
    28.59819, 25.8653,
  124.686, 125.2798, 123.8336, 120.9833, 117.8752, 115.3924, 114.5734,
    114.5908, 105.4935, 109.7312, 114.0058, 112.9368, 116.0212, 117.3371,
    107.4387, 87.779, 86.45618, 91.2361, 95.51884, 89.91563, 74.28064,
    58.96245, 54.47656, 41.64247, 34.17296, 31.2071, 28.09964, 27.1503,
    27.03773, 25.56988,
  110.1278, 100.569, 100.4526, 101.6036, 106.0853, 114.1703, 118.7743,
    119.4552, 116.3317, 116.9477, 116.0969, 115.7014, 117.0322, 117.1536,
    115.3574, 114.0699, 103.8036, 101.6505, 99.57731, 87.23225, 57.54195,
    50.86947, 39.48656, 33.2642, 30.89455, 29.60561, 27.36349, 25.81336,
    24.89169, 24.02316,
  95.03043, 97.61494, 102.4026, 106.2837, 110.4822, 117.3682, 120.2134,
    118.1633, 113.4887, 111.4661, 111.1989, 103.3707, 100.8465, 113.5577,
    109.1438, 103.795, 99.54542, 84.98375, 75.46453, 63.19958, 41.34293,
    39.76013, 33.30238, 31.89713, 30.78628, 28.75275, 26.70692, 25.68641,
    24.59758, 23.74816,
  85.22855, 84.25627, 87.62669, 92.13769, 95.82034, 100.0173, 102.9652,
    103.4456, 99.72795, 98.15236, 92.03152, 103.0738, 117.5659, 107.9495,
    100.9665, 91.39814, 80.56343, 67.54593, 63.50462, 57.20539, 36.49533,
    37.9996, 33.97921, 32.02603, 30.22931, 28.91217, 26.44178, 24.56373,
    24.05077, 23.64342,
  69.79138, 73.49062, 73.65903, 77.45045, 80.56109, 84.79814, 87.87971,
    89.76082, 92.07355, 92.79446, 106.8131, 119.5753, 119.4085, 117.4687,
    109.4938, 88.15517, 65.68685, 57.26422, 62.78687, 56.41794, 37.84219,
    38.95253, 34.97226, 32.84776, 29.09696, 27.51202, 26.10299, 23.68999,
    23.48731, 23.22716,
  76.78959, 74.39864, 65.17384, 62.61199, 66.22383, 69.60173, 74.37432,
    80.32506, 84.89783, 94.18749, 109.0452, 108.5528, 90.33266, 89.33363,
    83.03696, 74.84262, 75.71313, 79.77718, 81.37703, 68.16425, 47.49594,
    40.87726, 35.48365, 32.04198, 27.72413, 26.08124, 25.18566, 23.7004,
    23.30543, 23.15386,
  73.19768, 66.71243, 57.24107, 51.77594, 56.28989, 61.30872, 68.20998,
    75.31396, 83.47004, 95.55809, 97.50023, 77.10019, 69.856, 68.57118,
    65.75524, 66.77367, 73.25769, 80.15891, 79.07196, 72.40237, 58.40126,
    45.79129, 36.35077, 32.27212, 29.0357, 26.26686, 25.10631, 23.91173,
    23.27945, 23.17965,
  64.01833, 57.8484, 49.80824, 47.07776, 52.34921, 58.70929, 64.9389,
    70.83077, 77.16923, 82.35349, 73.49339, 57.72774, 63.7426, 64.37003,
    63.81768, 63.82076, 65.61006, 65.6218, 64.11418, 60.18701, 54.58964,
    50.63177, 42.4155, 35.89174, 31.33906, 27.77671, 25.16974, 23.99946,
    23.29696, 23.21345,
  63.22781, 53.58516, 49.04984, 48.95898, 54.10961, 56.20158, 61.61592,
    64.76074, 70.39044, 71.16759, 58.68987, 52.41263, 59.76522, 60.955,
    60.18662, 58.90971, 56.00278, 52.74141, 51.49619, 49.97372, 49.06945,
    47.9138, 45.95386, 44.2335, 37.37376, 29.23219, 25.39111, 24.40276,
    23.38148, 23.19315,
  60.43184, 55.043, 49.27926, 50.43616, 59.08699, 63.08744, 63.90631,
    60.45033, 61.75558, 58.94557, 47.50772, 50.33112, 54.91683, 56.24593,
    54.11841, 53.14362, 50.71202, 45.64177, 44.07775, 43.9597, 44.15414,
    43.57864, 41.64835, 42.50409, 41.31311, 32.84121, 26.89963, 26.57828,
    24.71722, 23.3378,
  63.97468, 61.39519, 62.3578, 65.98841, 71.17022, 70.85459, 71.29613,
    67.79836, 67.29015, 57.51637, 46.87871, 54.16505, 57.6778, 59.41843,
    56.79298, 54.72284, 52.65361, 48.12043, 43.78685, 42.90385, 42.08585,
    40.45924, 38.8864, 38.41335, 39.49417, 38.99151, 33.59691, 28.21718,
    26.31498, 24.12166,
  67.42169, 71.12029, 66.92783, 69.16679, 72.50784, 70.32523, 67.22453,
    66.79741, 70.4245, 61.20321, 48.84676, 56.25568, 59.21747, 61.24109,
    58.84883, 57.36395, 53.45226, 49.57349, 45.28821, 41.56629, 41.38671,
    41.22791, 38.74895, 36.34805, 36.12612, 39.40867, 39.44681, 33.31158,
    30.1142, 26.86694,
  79.58929, 84.74937, 82.92046, 77.51779, 72.5162, 69.17351, 72.63898,
    76.57919, 70.87579, 59.2726, 55.49828, 60.68931, 63.17349, 61.48737,
    56.73164, 55.09504, 52.45603, 49.34413, 46.73237, 43.02673, 42.46381,
    41.33053, 37.19278, 34.57556, 35.55799, 38.3339, 40.96457, 37.22413,
    29.95612, 26.62889,
  91.00816, 91.90907, 80.6827, 73.51822, 70.62318, 67.46038, 75.15739,
    75.101, 63.78553, 56.42835, 60.41551, 62.75861, 62.38385, 58.79942,
    55.22111, 53.06348, 50.26208, 47.578, 45.13571, 42.08518, 43.51721,
    46.71664, 46.2163, 43.32531, 43.36667, 45.17655, 48.15417, 44.02349,
    30.44968, 24.17888,
  93.06229, 86.88593, 77.1656, 75.84798, 76.29797, 74.43518, 76.27209,
    70.22742, 57.64765, 59.42533, 61.76457, 61.78932, 60.70707, 57.68087,
    55.96737, 52.59181, 48.15482, 46.92629, 48.69183, 51.35786, 53.84396,
    53.70686, 49.92763, 47.75166, 47.58964, 49.15962, 49.77416, 50.81796,
    43.18469, 27.64402,
  77.71059, 72.78047, 77.67885, 86.02945, 86.86415, 87.14418, 79.30347,
    63.03606, 54.90265, 56.44305, 52.59699, 50.94506, 51.60684, 52.68908,
    54.58022, 55.38359, 55.54364, 57.01607, 55.99928, 53.14571, 52.30417,
    49.28899, 45.25547, 43.24868, 44.06611, 45.22335, 44.60687, 42.04604,
    39.06444, 31.13577,
  76.70753, 79.25574, 81.36298, 81.09172, 82.52655, 88.57777, 85.53975,
    64.67831, 53.50798, 57.01535, 58.65237, 62.38773, 65.21129, 65.36787,
    63.90236, 62.56515, 57.68023, 51.79532, 48.71546, 45.15542, 42.03912,
    40.25018, 38.77163, 37.80195, 37.77349, 38.15269, 36.96185, 32.76433,
    28.72102, 24.38058,
  29.19157, 29.69408, 30.45255, 31.37376, 32.13591, 33.24316, 34.56416,
    35.97219, 37.58689, 39.67117, 42.63348, 43.81018, 41.83884, 43.23547,
    44.14277, 43.64664, 43.98324, 44.99178, 46.09612, 47.9488, 48.77754,
    47.44333, 48.19971, 50.60981, 51.98546, 51.34018, 54.86509, 55.55169,
    39.94102, 34.69554,
  31.15413, 32.38824, 32.88066, 35.04161, 35.92683, 37.24483, 39.41438,
    41.5396, 43.88259, 46.5085, 49.66986, 53.31219, 55.77235, 54.8205,
    54.31741, 55.11834, 54.37488, 55.87343, 57.78818, 59.54486, 59.85246,
    59.3209, 59.43336, 62.27158, 65.02036, 59.14378, 51.5262, 54.21523,
    40.69309, 36.09524,
  33.64194, 35.71684, 37.7663, 39.83067, 41.68473, 43.54056, 45.23484,
    47.05145, 49.00258, 50.94899, 53.05505, 55.73104, 58.40413, 61.12809,
    62.56805, 60.9423, 62.31424, 65.09045, 67.80338, 72.33412, 79.05877,
    84.45428, 84.03159, 80.15295, 76.37799, 70.88504, 62.43588, 51.51189,
    39.83282, 36.85569,
  40.55959, 43.45001, 46.64916, 49.73528, 52.26203, 54.63224, 55.55869,
    55.78551, 57.03739, 58.28036, 58.77745, 59.64172, 59.85789, 59.95202,
    63.81438, 65.83405, 63.40354, 62.15259, 67.16588, 73.09815, 81.36487,
    82.34256, 77.79915, 82.40472, 80.42995, 77.9391, 73.31926, 57.96827,
    43.45424, 35.65814,
  49.34086, 51.55305, 55.08537, 57.77422, 59.55292, 60.48692, 61.77589,
    62.98499, 65.48286, 67.36347, 67.73939, 70.21824, 71.79967, 72.12697,
    72.89662, 73.30536, 69.91691, 65.17085, 66.90167, 73.11035, 73.17473,
    64.44397, 66.52729, 73.15348, 79.10321, 79.68367, 75.6089, 80.36225,
    70.00296, 43.72736,
  62.26498, 67.40776, 71.68365, 75.55722, 74.84109, 74.08515, 77.01208,
    77.63292, 77.36938, 79.27716, 83.43658, 92.77125, 101.5992, 98.93785,
    98.94808, 99.24464, 96.12068, 86.53576, 75.12906, 72.48405, 64.40546,
    57.38339, 62.58442, 67.25347, 72.35735, 72.28086, 71.91031, 84.12207,
    73.37617, 39.44788,
  65.85649, 70.19159, 74.32335, 78.35236, 79.55469, 81.93799, 88.2087,
    92.86127, 91.11809, 86.22176, 82.20496, 73.35254, 63.82082, 65.71975,
    67.88089, 70.55044, 71.49129, 67.55699, 61.74619, 62.53059, 60.05692,
    59.5324, 63.41596, 68.82231, 69.17924, 64.36971, 67.76958, 74.46712,
    60.66338, 33.12705,
  59.68178, 63.84983, 68.96092, 73.75609, 76.02889, 82.84107, 85.70861,
    71.21427, 64.38976, 66.15529, 64.62923, 63.21495, 62.66645, 64.8604,
    66.54326, 68.95168, 71.39997, 69.62791, 64.68037, 64.55771, 64.94199,
    67.60005, 72.17096, 74.21017, 70.27007, 69.30363, 75.25264, 71.21674,
    51.61243, 34.63175,
  73.44775, 76.95745, 80.63628, 83.57969, 85.59185, 88.04732, 80.78915,
    82.12042, 87.31633, 90.11403, 91.07434, 91.36569, 93.49503, 101.5788,
    103.5609, 90.1954, 87.97459, 89.00945, 85.7547, 77.95488, 74.84048,
    81.23466, 87.68356, 84.54404, 75.83585, 79.97418, 77.83913, 61.92532,
    37.70586, 34.34067,
  102.821, 108.6472, 101.9941, 102.9917, 104.7976, 97.67093, 82.34708,
    90.34701, 91.32158, 95.38593, 99.61541, 104.6979, 102.1516, 97.79573,
    92.9373, 96.64854, 96.7115, 92.86417, 88.11151, 86.49687, 88.16982,
    83.42689, 76.81769, 68.60566, 72.93812, 80.4729, 69.16397, 44.67415,
    33.95801, 32.06046,
  116.9702, 115.9825, 117.0532, 111.0119, 116.1664, 110.0285, 101.3635,
    102.3845, 102.6198, 96.32007, 81.34314, 64.76572, 62.22594, 62.68185,
    63.22688, 65.2406, 67.98608, 68.92236, 69.27869, 72.93121, 81.40047,
    75.57629, 61.42745, 58.16847, 62.53046, 59.38593, 44.08865, 34.91717,
    34.46245, 32.21846,
  122.6944, 118.8983, 121.2999, 121.2385, 120.2075, 104.1864, 99.17844,
    90.05713, 80.87444, 71.60954, 66.31404, 63.31389, 65.94917, 66.5014,
    63.53472, 61.8973, 60.44631, 60.84612, 61.84341, 66.33054, 74.34573,
    71.39268, 60.68127, 68.01602, 68.86435, 52.6215, 36.4361, 39.44944,
    35.97215, 33.50349,
  127.9947, 127.8284, 129.1935, 129.3898, 127.8057, 123.6675, 116.4437,
    110.9421, 113.8377, 97.40526, 91.72336, 86.07165, 91.6034, 92.75487,
    81.46651, 67.63318, 68.43612, 66.78192, 65.92909, 69.90637, 71.30824,
    64.19924, 57.38536, 53.10618, 51.65529, 45.39545, 37.54432, 38.71306,
    37.92498, 34.82975,
  116.8432, 117.497, 117.7197, 117.3184, 117.009, 117.4931, 118.288,
    118.0791, 115.8575, 115.7377, 116.1537, 114.7449, 115.5221, 115.6667,
    106.5411, 85.71021, 80.34338, 83.49516, 84.67218, 76.42233, 64.54436,
    55.63341, 50.17459, 41.89676, 37.99181, 37.47166, 35.44117, 34.54673,
    34.97878, 34.04894,
  104.4229, 102.9596, 107.722, 111.1508, 114.075, 116.7721, 118.4281,
    117.7411, 110.7778, 108.1371, 100.9195, 94.50639, 95.95544, 98.23689,
    95.763, 91.74116, 81.09531, 76.69456, 75.394, 68.09177, 52.27453,
    50.23835, 43.05125, 40.10206, 38.97332, 37.40515, 35.75439, 34.32784,
    33.35319, 32.75619,
  103.3821, 107.8873, 109.5005, 109.6022, 107.6828, 107.5399, 108.6314,
    99.98491, 88.61832, 83.34864, 81.44244, 75.6906, 72.63896, 79.21028,
    76.1599, 73.06387, 72.87285, 65.5454, 62.36172, 55.72092, 44.63884,
    45.76998, 41.29746, 39.78459, 38.97919, 37.27027, 35.42929, 34.54864,
    33.58166, 32.77832,
  86.78671, 86.12915, 88.33176, 90.27312, 91.61317, 93.25828, 93.39763,
    92.4792, 88.88264, 83.69407, 76.84624, 84.24519, 91.05184, 82.40449,
    75.74072, 69.6722, 64.17793, 60.41001, 60.80494, 55.74237, 44.34104,
    45.67411, 42.04561, 39.68261, 38.37939, 37.24089, 34.74531, 33.05355,
    32.92899, 32.61548,
  79.17536, 82.13226, 81.08849, 82.7413, 83.81622, 85.25774, 85.63994,
    85.7453, 87.79477, 87.99916, 96.9275, 104.5868, 100.2586, 96.37073,
    90.21954, 78.90143, 68.57695, 66.22296, 67.9912, 59.96386, 45.57779,
    44.75708, 41.99529, 40.25599, 37.0803, 35.70963, 34.68308, 32.5596,
    32.46449, 32.27155,
  89.28739, 81.99516, 69.94139, 64.00502, 64.46902, 64.39143, 66.19561,
    69.08455, 70.77394, 75.98215, 82.8474, 81.16689, 73.28639, 77.74107,
    79.33812, 82.03076, 88.02612, 92.43195, 88.73672, 76.1408, 56.99025,
    48.21235, 43.53098, 40.46704, 37.08437, 35.19432, 34.27768, 32.93661,
    32.45834, 32.29384,
  81.34824, 73.6951, 62.9631, 56.35652, 58.67968, 60.69893, 63.4053,
    65.78404, 69.37021, 75.35625, 74.1414, 63.09774, 62.77241, 62.3409,
    61.93233, 62.41512, 67.30318, 73.59548, 75.9207, 74.05782, 65.86526,
    55.69577, 47.10836, 43.05857, 39.63597, 36.03718, 34.46358, 33.12677,
    32.45557, 32.31654,
  75.42635, 67.78807, 58.61213, 54.59407, 56.54416, 58.16965, 59.18038,
    60.09415, 62.10174, 63.51252, 57.92174, 50.35788, 54.81419, 54.36192,
    52.64044, 51.75898, 53.35422, 56.06599, 59.5192, 61.21668, 61.53228,
    60.96898, 54.75053, 48.01714, 42.42893, 37.34563, 34.45306, 33.19173,
    32.45728, 32.3298,
  76.45441, 68.53238, 61.32212, 58.27045, 58.99026, 56.39774, 56.29077,
    55.62083, 57.8848, 57.01133, 48.30565, 44.36786, 47.25031, 47.47497,
    46.67677, 47.07023, 47.1082, 48.32682, 51.12398, 53.14948, 54.20751,
    54.3462, 55.15752, 54.21316, 47.55572, 38.98177, 35.27401, 34.13055,
    32.72911, 32.29901,
  80.12508, 76.18217, 66.90839, 64.27107, 66.8095, 65.57544, 62.46443,
    57.06588, 56.9837, 53.79358, 46.51896, 47.46457, 48.93105, 49.57769,
    48.74725, 49.82877, 49.82918, 47.63116, 47.8697, 48.92686, 49.58944,
    49.80394, 49.66345, 51.79688, 52.20372, 44.61125, 38.18305, 36.64441,
    34.40676, 32.48944,
  88.43878, 85.65984, 80.77774, 78.92252, 78.92252, 76.86091, 75.94846,
    74.83636, 73.99925, 66.38105, 58.78807, 62.89391, 64.32054, 65.4472,
    63.2991, 61.84088, 60.328, 56.80228, 53.15728, 52.23007, 51.37532,
    50.52796, 49.86407, 49.67588, 51.69723, 52.04758, 46.07574, 39.34905,
    36.89188, 33.6961,
  85.45294, 82.58975, 73.73776, 71.94017, 72.1512, 70.87955, 71.40112,
    73.95178, 77.70466, 69.15727, 61.02539, 64.74611, 67.08379, 68.14967,
    66.70692, 65.68769, 62.83513, 60.49694, 58.28031, 55.77037, 54.31936,
    52.43115, 49.46725, 47.78252, 48.93339, 51.9697, 51.86596, 44.45044,
    39.62744, 35.84273,
  93.27442, 89.73169, 83.4563, 76.91298, 73.25481, 72.22711, 76.7115,
    79.97977, 75.61185, 67.42358, 66.39523, 68.33707, 70.25165, 69.05303,
    66.34705, 65.7468, 64.52757, 63.25516, 63.15044, 61.7543, 60.25289,
    58.09531, 53.94758, 50.93621, 51.43655, 52.75288, 53.46054, 46.33735,
    37.43902, 34.66179,
  94.58181, 89.27666, 80.31522, 75.5136, 72.08325, 68.49698, 72.8991,
    73.44244, 68.36835, 65.39418, 69.06863, 71.29082, 72.35939, 71.87032,
    70.41872, 69.04768, 67.35855, 67.07807, 67.61407, 67.11273, 67.14053,
    68.06378, 66.66481, 63.20861, 62.63149, 63.60912, 64.62115, 56.88517,
    40.88572, 33.03537,
  93.80313, 88.21051, 84.28406, 82.83537, 80.49532, 76.67346, 74.69956,
    70.38931, 64.06893, 66.57658, 68.90306, 71.11589, 72.08089, 71.72615,
    71.32565, 69.21624, 65.92948, 64.97421, 66.22041, 66.7336, 63.69537,
    59.59827, 56.27956, 55.47902, 56.8007, 58.41415, 59.38969, 60.78638,
    52.88739, 36.97874,
  79.42493, 77.2121, 80.05479, 83.31711, 85.89366, 86.85548, 79.12967,
    66.72365, 61.92475, 62.40815, 60.26786, 59.57413, 59.87475, 59.94456,
    59.88974, 59.19948, 56.81452, 54.74478, 52.05906, 48.84314, 47.52647,
    46.09071, 43.59563, 42.10115, 43.23437, 44.46593, 44.29486, 42.76001,
    42.84823, 38.25581,
  68.63759, 70.19568, 70.07832, 69.73337, 74.28787, 81.36122, 80.6464,
    65.85608, 58.6461, 61.76122, 62.88713, 63.79602, 63.13579, 59.96267,
    55.98548, 52.46301, 46.48937, 41.32299, 40.53921, 39.58475, 37.95226,
    38.26656, 38.27585, 38.16991, 38.62669, 39.75061, 39.69845, 37.19135,
    34.47145, 32.29131,
  42.05692, 42.89197, 43.51875, 44.20557, 44.62959, 45.16499, 45.77893,
    46.39731, 47.12351, 48.01243, 49.32468, 49.32226, 47.13032, 47.35617,
    47.3022, 46.49451, 46.32407, 46.7299, 47.27714, 48.18881, 48.24252,
    46.82567, 47.2301, 49.12324, 50.37256, 49.595, 51.66254, 52.81171,
    42.12257, 38.35085,
  47.83998, 48.92273, 48.97118, 50.16459, 50.29876, 50.6689, 51.63976,
    52.57964, 53.5785, 54.68481, 55.94616, 57.42331, 58.17145, 56.80111,
    55.89096, 56.04624, 55.18121, 56.00127, 57.17038, 58.08609, 57.74562,
    56.77118, 56.5801, 58.76448, 61.12063, 55.90194, 48.62783, 51.44622,
    42.49456, 39.21138,
  50.19081, 51.23082, 51.82026, 52.39258, 52.87219, 53.44356, 54.02234,
    54.78796, 55.59101, 56.36572, 57.28545, 58.61915, 59.92874, 61.45153,
    62.17683, 60.86267, 61.56596, 63.47258, 65.50791, 68.54113, 73.35911,
    77.45214, 76.85828, 73.12112, 69.5535, 64.78513, 57.91038, 49.60299,
    41.91327, 39.88066,
  55.2844, 56.35488, 57.40371, 58.47451, 59.17142, 59.96786, 59.98979,
    59.63103, 59.93559, 60.23307, 60.15137, 60.40031, 60.1396, 59.726,
    62.01875, 63.17748, 61.32873, 60.72919, 64.34201, 68.32211, 74.35528,
    74.75549, 69.93256, 73.01746, 70.92795, 69.30389, 66.7654, 55.39532,
    44.52926, 39.04136,
  61.66923, 61.84361, 63.06699, 63.81112, 63.91632, 63.89963, 64.34518,
    64.63243, 65.76128, 66.53139, 66.69798, 68.42372, 69.06595, 68.52211,
    68.74221, 69.30688, 66.81615, 63.199, 64.15634, 68.49106, 68.22812,
    60.40004, 61.49207, 66.45892, 70.89521, 71.6935, 69.86887, 74.71384,
    67.63138, 46.17123,
  66.03555, 68.63216, 70.91119, 72.9372, 71.97104, 71.56116, 73.96504,
    74.46114, 73.78812, 74.61055, 77.7241, 85.45724, 92.3671, 89.10135,
    89.1881, 90.0706, 87.4179, 79.93457, 71.12962, 68.3675, 61.17937,
    54.73425, 58.55286, 61.8991, 65.92791, 66.85835, 67.74979, 77.71499,
    70.20912, 42.70098,
  68.33215, 71.82962, 74.61792, 77.21051, 77.92461, 80.23991, 86.16208,
    90.51633, 88.88464, 84.16653, 80.1713, 71.93361, 62.56436, 63.01785,
    64.12257, 66.21906, 66.89497, 63.97344, 59.76847, 59.79955, 57.34736,
    56.24324, 58.70063, 62.44712, 63.0752, 60.2574, 63.55652, 70.28378,
    59.7081, 37.06519,
  73.48512, 76.71854, 79.53545, 82.1076, 82.981, 87.75305, 89.55663,
    76.48816, 69.69126, 69.7194, 67.05559, 64.12552, 61.97654, 61.93184,
    61.96127, 63.34615, 65.62906, 64.61824, 61.21984, 60.44783, 60.2373,
    61.78948, 64.74036, 66.32623, 64.08794, 63.91666, 69.07738, 66.93845,
    51.07982, 37.95501,
  82.18246, 83.12395, 83.66239, 84.1349, 84.94699, 85.3343, 76.89254,
    75.94644, 78.13795, 78.11119, 77.82751, 77.13295, 77.46518, 82.23029,
    83.68742, 75.584, 75.05792, 76.4798, 74.53724, 69.03167, 66.13017,
    69.74514, 74.08498, 72.31302, 67.38692, 71.43605, 71.02347, 59.39796,
    40.03048, 38.06788,
  94.81862, 96.07367, 89.07648, 88.11247, 87.64484, 81.45138, 66.9287,
    71.98657, 71.22647, 72.50748, 74.12565, 77.58492, 77.16846, 75.74062,
    74.22415, 77.96219, 79.00698, 77.39303, 74.86271, 73.68671, 74.42798,
    71.02223, 66.69794, 62.04726, 65.86171, 73.20793, 66.10773, 45.56672,
    37.72643, 36.56317,
  113.5393, 112.8182, 112.0825, 98.78658, 98.49718, 89.02392, 80.32816,
    80.76578, 81.3455, 77.6311, 67.78046, 56.71096, 55.39972, 56.33027,
    57.36881, 59.02081, 61.08083, 62.06701, 62.81099, 65.23744, 70.8665,
    67.35832, 58.3194, 57.04018, 60.88813, 58.74038, 45.99226, 38.15991,
    38.12804, 36.64588,
  121.3051, 118.1853, 119.6649, 118.5358, 115.8609, 97.70747, 91.17789,
    82.50367, 75.8231, 70.40805, 65.52392, 62.6088, 63.99688, 63.3577,
    59.48986, 58.51344, 57.51337, 57.4938, 57.93484, 60.87608, 66.21862,
    64.54636, 57.87606, 63.98129, 65.79408, 52.90254, 39.4421, 41.74888,
    39.0432, 37.4765,
  123.1557, 123.4016, 123.9445, 123.4916, 121.3493, 117.5512, 111.1831,
    101.104, 103.7881, 91.89993, 86.11221, 80.73656, 84.80609, 84.92813,
    75.52721, 63.29839, 63.9852, 62.7999, 61.45292, 63.05238, 63.90459,
    59.83355, 55.64042, 51.8794, 50.85807, 46.62879, 40.43096, 41.22212,
    40.55558, 38.43871,
  109.8297, 110.3441, 107.1834, 104.1283, 103.2534, 109.7784, 111.8822,
    111.4435, 101.7201, 102.4194, 106.928, 102.0316, 100.9413, 100.1332,
    91.38185, 77.24756, 71.27957, 75.08981, 76.21652, 69.20336, 60.56931,
    54.23165, 49.6078, 43.30165, 40.33546, 40.19076, 38.99201, 38.2923,
    38.56171, 37.8947,
  78.07925, 75.14943, 76.68048, 77.45461, 78.6936, 80.48909, 85.61269,
    85.71797, 81.09741, 81.35341, 77.50224, 75.03207, 77.67276, 80.97047,
    80.37752, 78.43913, 72.25263, 68.45924, 67.05601, 62.12383, 51.27896,
    49.73993, 43.99709, 41.68563, 41.07069, 40.24791, 39.13451, 38.09789,
    37.38339, 36.94736,
  76.66924, 78.70493, 78.96208, 78.38297, 77.63609, 79.40707, 81.49365,
    77.02042, 71.93865, 68.97374, 68.24303, 65.06501, 63.82104, 67.9696,
    65.69833, 64.4602, 64.78195, 59.72001, 56.88116, 52.46933, 45.19869,
    45.54021, 42.36929, 41.34174, 41.04868, 40.1786, 38.95994, 38.21095,
    37.51368, 36.9736,
  69.32494, 68.62704, 69.41636, 71.10958, 72.65854, 74.11569, 76.17076,
    78.22163, 76.37102, 72.93076, 68.88638, 73.85368, 78.27454, 73.2114,
    67.36191, 63.0542, 59.44271, 56.78623, 55.75548, 52.45443, 45.31274,
    45.66929, 42.86158, 41.30401, 40.62943, 40.1238, 38.50358, 37.23487,
    37.09967, 36.87463,
  64.78217, 65.50311, 64.56381, 66.47161, 68.41563, 70.95965, 73.02498,
    75.03462, 76.29514, 75.73518, 80.5421, 84.65322, 83.22315, 82.29239,
    77.98132, 72.40494, 66.83922, 64.62771, 63.68698, 56.93727, 46.77974,
    45.16161, 43.02009, 41.9239, 40.01224, 39.15677, 38.37734, 36.89663,
    36.7782, 36.65276,
  71.41075, 66.12578, 58.62984, 55.38419, 57.71346, 58.67047, 60.47041,
    62.19894, 62.73245, 65.23875, 69.06465, 67.78638, 63.53744, 66.36056,
    67.89014, 70.51885, 76.39482, 80.39075, 77.75876, 68.70738, 55.50472,
    47.99866, 44.19664, 42.45416, 40.25125, 38.92316, 38.1759, 37.10566,
    36.76929, 36.68395,
  64.89488, 59.87984, 52.80744, 48.69574, 50.45423, 51.45904, 52.9097,
    54.47867, 56.88934, 60.92129, 60.98625, 55.38723, 55.75858, 55.24121,
    54.72677, 55.34903, 59.14537, 64.34218, 66.27469, 65.15286, 59.78593,
    52.76672, 46.84367, 44.26199, 41.98791, 39.55906, 38.35441, 37.28357,
    36.76396, 36.67935,
  61.83983, 57.34084, 50.23628, 46.65412, 47.57701, 48.33288, 49.54068,
    51.0214, 53.29883, 55.39819, 52.74242, 49.31171, 52.23083, 52.0472,
    50.78225, 50.31251, 51.5979, 53.42295, 55.25335, 55.35247, 55.02289,
    54.83926, 51.49597, 47.45417, 43.87649, 40.47013, 38.37355, 37.31954,
    36.76148, 36.69002,
  66.54501, 62.70269, 55.5183, 52.60408, 52.93135, 51.50426, 51.85976,
    52.22201, 54.67386, 54.98429, 50.25927, 47.89268, 49.58625, 49.58591,
    49.02616, 49.11354, 48.90062, 49.32432, 50.61696, 51.15757, 51.04893,
    50.78986, 51.22136, 50.88682, 46.88823, 41.46466, 38.94576, 37.94524,
    36.93459, 36.65598,
  74.14249, 73.55714, 65.23782, 63.14277, 65.20851, 64.87628, 62.48175,
    59.74802, 59.80927, 57.83545, 53.29381, 53.67929, 54.02795, 53.89074,
    52.70226, 52.73446, 52.07867, 50.04198, 49.51641, 49.31421, 48.72342,
    48.22601, 47.91403, 49.03704, 49.51259, 44.97486, 40.87062, 39.62126,
    38.03096, 36.77803,
  79.46862, 78.97797, 74.15323, 72.68529, 72.8655, 71.65348, 71.75526,
    71.18261, 72.5359, 68.06525, 63.20856, 65.00928, 65.86018, 65.72829,
    63.69655, 62.05194, 59.97551, 56.95712, 53.78697, 52.01126, 50.38615,
    49.12438, 48.23053, 47.97912, 49.24789, 49.69041, 46.12865, 41.48181,
    39.72111, 37.57681,
  80.7991, 76.73241, 70.19899, 68.21143, 68.48476, 68.11189, 69.11993,
    72.31404, 76.00182, 71.10526, 65.16629, 66.91973, 67.70834, 67.8428,
    66.48257, 65.23888, 62.49094, 59.97484, 57.53123, 54.76888, 52.92402,
    50.95339, 48.33379, 46.81328, 47.64325, 49.73012, 49.86218, 44.95589,
    41.52176, 38.96172,
  85.70056, 82.78365, 77.4272, 72.3001, 69.8116, 68.97691, 72.62285,
    76.75121, 75.68893, 70.49684, 69.38321, 69.90706, 70.24243, 68.84527,
    66.67216, 65.742, 64.26991, 62.55561, 61.09945, 58.80687, 57.46732,
    55.73944, 51.94885, 49.26213, 49.3289, 50.15262, 50.73314, 46.27071,
    40.2354, 38.19398,
  85.17126, 81.62434, 75.19362, 71.01573, 67.89407, 65.05185, 68.20175,
    69.38595, 67.08945, 65.07126, 66.73888, 67.82489, 68.27004, 67.70501,
    66.51955, 65.28352, 63.96262, 63.16432, 62.29322, 61.00969, 61.00379,
    61.66159, 59.94493, 56.789, 56.0192, 56.73854, 57.47957, 52.63712,
    42.29186, 37.17509,
  78.08064, 75.51262, 72.04427, 70.56435, 69.79885, 66.03073, 63.71299,
    60.50252, 56.72284, 57.3163, 58.39629, 59.97466, 61.37287, 62.07943,
    62.2969, 61.4307, 59.79851, 59.18747, 59.60331, 59.68805, 58.30651,
    55.91808, 53.04827, 51.9398, 52.62077, 53.75329, 54.16872, 54.8938,
    49.7536, 39.70766,
  61.48642, 61.24228, 62.43321, 63.407, 65.58805, 67.01988, 61.68702,
    53.2678, 50.64563, 51.62638, 51.27361, 51.50843, 52.32875, 52.89737,
    53.29397, 53.30099, 52.31922, 51.51815, 49.96357, 48.13282, 47.48115,
    46.63458, 45.01318, 43.99136, 44.81411, 45.47198, 44.97163, 43.67385,
    43.51922, 40.53991,
  51.15804, 51.72127, 51.48838, 50.75318, 53.24703, 58.0312, 58.34062,
    50.46154, 46.80691, 49.37844, 51.20998, 52.70832, 52.94267, 51.49949,
    49.55383, 48.18161, 45.19817, 42.35237, 42.03013, 41.41938, 40.49318,
    40.88306, 41.11194, 41.15809, 41.39073, 41.91988, 41.60428, 39.97226,
    38.25707, 36.74791,
  40.84348, 41.08062, 41.25468, 41.46924, 41.59064, 41.77989, 42.05637,
    42.32446, 42.69666, 43.42013, 44.49419, 44.26128, 42.40236, 42.93062,
    43.16658, 42.78145, 43.00912, 43.57352, 44.23377, 45.35184, 45.83521,
    44.98725, 45.5602, 47.3691, 48.85846, 48.80648, 50.54645, 51.37041,
    43.27151, 40.36037,
  45.39079, 45.71083, 45.27659, 45.78957, 45.53182, 45.42928, 45.66737,
    45.81881, 46.15969, 46.70051, 47.42675, 48.23654, 48.59826, 47.54031,
    46.9409, 47.4602, 47.09385, 47.96207, 49.07233, 50.03635, 50.35204,
    50.50733, 51.78852, 55.25872, 58.22406, 54.10728, 47.93848, 50.74528,
    43.57903, 40.98703,
  48.2485, 48.64701, 48.7745, 48.9579, 49.15195, 49.43064, 49.67003,
    50.01231, 50.51426, 51.13725, 51.80267, 52.82126, 53.9618, 55.34624,
    56.14627, 55.43155, 56.374, 58.04287, 59.57105, 62.15542, 66.85921,
    71.67458, 72.14407, 68.84557, 65.81381, 61.60625, 55.93064, 49.79118,
    43.47292, 41.75033,
  52.19135, 52.94498, 53.73761, 54.60217, 55.22831, 56.06548, 56.1652,
    55.9371, 56.40064, 56.95708, 57.22511, 58.01035, 58.29638, 58.11062,
    60.29655, 61.46022, 60.18434, 59.80684, 62.7201, 66.27461, 71.87346,
    71.81178, 66.43559, 68.00271, 64.98139, 63.38423, 62.20334, 52.69108,
    44.0759, 40.6867,
  55.24823, 55.06879, 55.89831, 56.46616, 56.76726, 56.82551, 57.23792,
    57.5895, 58.63097, 59.15877, 59.05937, 60.48296, 61.40373, 61.66234,
    62.59447, 63.90708, 63.09497, 61.55341, 63.90496, 68.66818, 68.4015,
    60.36025, 60.1219, 64.12444, 66.99015, 67.08426, 65.5702, 70.06517,
    65.40469, 47.88352,
  61.46612, 63.6072, 65.61356, 67.60776, 67.41687, 67.83257, 70.4213,
    71.4628, 72.31989, 74.27574, 77.93472, 86.07525, 93.18564, 90.05397,
    90.05862, 90.95277, 88.41389, 81.2896, 73.07108, 70.26221, 63.50078,
    56.73113, 60.63503, 63.68092, 67.42126, 68.2533, 69.01617, 78.88552,
    72.41902, 44.85792,
  67.52962, 70.56437, 73.13666, 75.73131, 77.05707, 80.15955, 86.79798,
    91.93453, 91.01668, 86.67383, 82.89677, 75.32962, 66.76778, 67.43143,
    68.34058, 69.62911, 69.99438, 66.36979, 61.44482, 60.38177, 57.32677,
    56.19506, 58.9126, 62.52624, 63.74999, 62.05662, 65.76213, 71.79221,
    60.49377, 39.30417,
  66.16422, 68.41237, 70.68761, 73.02355, 74.01972, 78.56757, 80.37816,
    67.9324, 61.28048, 61.16304, 58.71064, 56.21306, 54.80233, 55.65578,
    56.89872, 59.25361, 61.74416, 61.32652, 58.40927, 57.90802, 57.51355,
    58.73144, 61.70366, 63.93607, 63.21484, 64.29992, 70.14111, 68.57635,
    53.0906, 39.62297,
  70.88102, 72.15629, 73.35216, 74.40439, 75.91022, 76.52209, 68.36896,
    66.7933, 68.63451, 68.73106, 68.72034, 68.59597, 69.57513, 74.04811,
    76.04977, 70.53841, 71.53533, 73.59348, 72.07018, 67.19681, 64.92885,
    68.25947, 72.05498, 70.77769, 67.29045, 71.9166, 72.87762, 61.43331,
    41.96849, 40.22529,
  82.55858, 85.98872, 81.6778, 82.57603, 84.32378, 79.08894, 66.48158,
    71.78742, 71.8615, 74.04823, 76.33807, 80.0451, 79.44105, 77.32001,
    75.15359, 77.68767, 78.32686, 76.90716, 74.65636, 73.85143, 74.29492,
    71.49043, 68.07256, 63.92344, 68.12828, 75.47009, 67.87084, 47.80688,
    39.63002, 38.96839,
  104.7702, 103.2153, 98.72552, 88.81902, 90.75249, 82.97707, 75.45688,
    77.85271, 78.95222, 76.41855, 68.67832, 59.07008, 58.22224, 58.96815,
    59.37064, 60.63552, 62.10298, 62.45357, 62.85316, 64.97421, 69.58044,
    66.39281, 58.72343, 57.68845, 62.15366, 60.97113, 48.49565, 39.70305,
    40.20935, 38.99248,
  109.9805, 107.1325, 109.1903, 108.7623, 101.3968, 83.22125, 80.35251,
    73.2676, 67.14407, 64.1887, 60.29193, 58.58512, 60.35524, 60.16919,
    58.01735, 57.90181, 57.37686, 57.74728, 58.25566, 60.83342, 65.82661,
    65.1124, 60.32641, 66.29836, 67.63936, 54.4052, 40.73923, 43.04022,
    40.80233, 39.63772,
  116.4651, 116.794, 117.5778, 116.747, 114.1248, 110.3485, 99.9374,
    84.41328, 90.13898, 79.49879, 75.27823, 71.68852, 75.71313, 76.6053,
    70.40667, 60.50071, 61.37572, 61.19885, 60.90211, 63.02706, 65.06908,
    62.88365, 59.57419, 56.62171, 54.65219, 48.94355, 42.33969, 43.32283,
    42.37125, 40.5652,
  107.5308, 107.8587, 107.4019, 105.4424, 103.9429, 103.7815, 104.0121,
    103.6373, 97.14442, 97.04317, 101.2933, 96.96547, 94.6152, 95.57299,
    87.75447, 73.81159, 70.71845, 73.65237, 75.39177, 68.83246, 61.16962,
    56.09256, 52.10606, 45.87959, 42.85634, 42.49471, 41.36893, 40.78585,
    40.85696, 40.17607,
  82.17524, 79.28851, 81.15061, 81.55646, 82.90139, 85.16054, 89.3028,
    88.46906, 84.08795, 84.30472, 80.85272, 77.4311, 79.49332, 82.66071,
    82.78296, 79.47311, 71.95174, 68.72438, 66.69405, 61.90635, 52.19707,
    50.23656, 45.22721, 42.96388, 42.6248, 42.03076, 41.17318, 40.31543,
    39.71398, 39.32218,
  73.26918, 75.48299, 76.00785, 75.51282, 74.48825, 75.50248, 77.00504,
    73.74915, 69.53777, 66.83922, 66.51212, 64.1275, 63.2804, 67.26688,
    65.36913, 63.75814, 63.96292, 59.131, 56.41923, 52.39558, 46.18487,
    46.45238, 43.73765, 42.75509, 42.58165, 42.01202, 41.13165, 40.41941,
    39.76105, 39.31161,
  64.77215, 63.84532, 64.26296, 65.29633, 66.24171, 66.87456, 68.03072,
    69.50403, 68.25412, 65.67108, 62.36922, 66.17184, 70.32597, 67.07605,
    62.87467, 60.21502, 57.67211, 55.65923, 54.93764, 52.34074, 46.22467,
    46.47748, 44.05569, 42.74731, 42.40558, 42.09464, 40.75375, 39.68131,
    39.46344, 39.23802,
  62.14401, 62.90191, 62.05485, 63.23787, 64.24245, 65.65651, 66.88041,
    68.345, 69.15077, 68.42125, 71.60513, 74.4359, 73.36704, 72.27676,
    68.04314, 63.53175, 59.02003, 57.81567, 58.32851, 53.9419, 46.63168,
    45.81915, 44.02157, 43.16016, 41.90285, 41.23486, 40.52303, 39.28776,
    39.1828, 39.06219,
  70.76875, 66.72939, 60.00359, 56.99449, 58.82673, 59.37882, 60.57312,
    61.80461, 62.09291, 64.0331, 67.18185, 66.19862, 62.26891, 63.79516,
    64.06315, 65.88198, 70.27424, 73.55034, 71.75884, 64.35959, 53.91914,
    47.91624, 44.779, 43.53699, 42.01692, 41.02164, 40.35372, 39.41737,
    39.13831, 39.07083,
  67.14194, 63.35072, 56.94992, 53.47543, 55.1585, 56.05867, 57.10434,
    58.08606, 59.90051, 63.28923, 63.5997, 59.09581, 59.04848, 58.23465,
    57.3583, 57.57464, 60.21177, 63.81296, 64.44253, 62.40858, 57.49708,
    51.4718, 46.69786, 44.99372, 43.47649, 41.54699, 40.5549, 39.5597,
    39.10337, 39.08181,
  63.43327, 59.86745, 53.39591, 50.18067, 51.08033, 51.66063, 52.45152,
    53.36345, 55.05183, 56.92664, 55.08745, 52.40129, 54.64574, 54.20758,
    53.02248, 52.46188, 53.09564, 54.05528, 54.8423, 54.23123, 53.60829,
    53.15034, 50.09667, 47.21469, 44.85004, 42.24978, 40.60042, 39.59666,
    39.11844, 39.07235,
  62.95417, 59.66281, 53.35077, 50.48629, 50.85757, 49.9619, 50.60421,
    51.04675, 53.0364, 53.44371, 50.03455, 48.53518, 50.07014, 50.18408,
    49.87213, 50.03569, 49.89869, 50.23033, 51.15924, 51.59204, 51.52869,
    51.16341, 51.03782, 49.95776, 46.76416, 42.87004, 41.0037, 40.0669,
    39.19281, 39.022,
  66.15619, 65.02727, 57.82701, 55.28568, 56.74626, 56.5463, 55.18944,
    53.31483, 53.51991, 52.25144, 49.05576, 49.59276, 50.28429, 50.61234,
    50.20291, 50.63678, 50.54219, 49.3546, 49.18356, 49.25924, 48.99166,
    48.62831, 48.04133, 48.42765, 48.46283, 45.11584, 42.32366, 41.30878,
    39.98391, 39.10821,
  72.56391, 72.1312, 67.28938, 65.27962, 65.00351, 63.52786, 63.57265,
    63.11195, 64.42186, 61.59281, 58.2633, 59.85442, 60.7255, 60.97025,
    59.68978, 58.56246, 57.33532, 55.13156, 52.68777, 51.35157, 50.25102,
    49.51051, 48.48843, 47.77602, 48.5767, 48.93785, 46.23854, 42.57937,
    41.18334, 39.71541,
  74.80544, 71.09779, 65.18589, 62.74174, 62.72234, 61.96328, 62.74677,
    65.51513, 68.65977, 65.13021, 60.8961, 62.49642, 63.62434, 64.15894,
    63.16774, 62.39897, 60.84119, 59.18736, 56.65816, 54.32249, 53.2037,
    51.83421, 49.35594, 47.78661, 48.50861, 50.31086, 50.12156, 45.67376,
    42.81177, 40.87431,
  77.85873, 75.09002, 70.17589, 65.36494, 63.77333, 63.11292, 65.91272,
    69.38576, 68.86871, 64.591, 63.80281, 64.45994, 65.19457, 64.47565,
    62.5752, 61.81679, 61.40747, 60.23511, 58.06631, 55.84468, 55.11221,
    54.04147, 50.87518, 48.82041, 49.15788, 49.92073, 50.44007, 46.77252,
    41.98555, 40.37957,
  79.03437, 75.51472, 70.26211, 66.48111, 64.71608, 63.15545, 66.22808,
    67.62955, 66.20772, 64.43096, 65.44341, 65.84857, 66.18631, 65.68971,
    64.34387, 63.43704, 63.09012, 62.48163, 60.62727, 59.15541, 59.81567,
    60.65079, 58.6301, 55.85423, 54.82991, 54.89237, 55.15505, 51.04202,
    42.94546, 39.42036,
  75.08849, 73.00281, 70.05156, 69.20664, 69.42844, 67.98763, 67.24467,
    65.2689, 62.53232, 63.10163, 63.99957, 65.0472, 66.02223, 66.51552,
    66.18797, 65.3131, 64.49371, 63.73249, 62.88546, 62.24173, 60.97837,
    58.80134, 56.0584, 54.6886, 54.64845, 54.57285, 54.12577, 53.89618,
    49.35486, 41.32729,
  62.65977, 62.84118, 63.71138, 64.60353, 66.5507, 68.15213, 64.47977,
    57.6719, 55.67948, 56.20662, 55.79966, 56.02618, 56.94575, 57.99705,
    58.60642, 58.67419, 57.84675, 56.70483, 54.48621, 52.03964, 50.79757,
    49.86079, 48.41437, 47.46568, 47.8676, 47.88968, 47.03748, 45.75051,
    45.18977, 42.44416,
  56.53633, 57.13331, 57.222, 56.93842, 59.12129, 63.28138, 63.21492,
    56.2084, 53.31853, 55.35556, 56.46823, 57.27252, 57.18449, 55.87606,
    54.08546, 52.69051, 49.81634, 47.23217, 46.60541, 45.49517, 44.36693,
    44.59483, 44.8096, 44.71012, 44.67476, 44.7043, 43.96468, 42.27418,
    40.71464, 39.22864,
  41.23412, 41.25696, 41.36527, 41.41862, 41.42308, 41.48349, 41.65042,
    41.90843, 42.23132, 42.74353, 43.58599, 43.45544, 42.00082, 42.3318,
    42.44382, 42.02829, 42.00564, 42.17224, 42.44882, 43.15898, 43.58017,
    43.10196, 43.55606, 45.07875, 46.66354, 47.03302, 48.65408, 50.06783,
    44.41794, 42.2032,
  42.33178, 42.45807, 42.1963, 42.58558, 42.37522, 42.28535, 42.58529,
    42.90569, 43.29898, 43.75647, 44.28214, 44.797, 44.97365, 44.08007,
    43.48672, 43.76621, 43.19931, 43.6825, 44.47895, 45.31347, 45.74189,
    46.4373, 48.49186, 53.08064, 57.23322, 53.57408, 47.98743, 50.70199,
    44.98663, 42.79533,
  42.16286, 42.13352, 42.18781, 42.29259, 42.3301, 42.4948, 42.73291,
    43.05135, 43.4219, 43.80189, 44.31918, 45.024, 45.73129, 46.66203,
    47.31269, 46.94307, 47.96975, 49.72241, 51.4329, 54.41052, 59.62981,
    65.80399, 68.11176, 66.86012, 64.9997, 59.8807, 55.08255, 50.02543,
    44.98803, 43.47844,
  43.57492, 44.11184, 44.93702, 45.82194, 46.57013, 47.39959, 47.62333,
    47.61502, 48.03876, 48.72432, 49.27468, 50.18738, 50.8998, 51.38073,
    53.86578, 55.83382, 55.88428, 56.593, 60.16323, 64.80675, 71.30778,
    71.84335, 66.20632, 66.91695, 63.73043, 61.64754, 60.08749, 51.94153,
    44.67667, 42.43828,
  47.41405, 47.57485, 48.62709, 49.38676, 49.7065, 49.65834, 49.668,
    49.56657, 50.03173, 50.22034, 50.13367, 51.47415, 52.88237, 54.46722,
    56.60909, 59.00746, 59.72781, 59.75479, 63.07184, 68.06485, 67.94565,
    59.60849, 57.59467, 61.12128, 63.36886, 63.18384, 62.40447, 67.30519,
    64.37937, 49.44198,
  48.80912, 49.69989, 51.02089, 52.18031, 51.6517, 51.45206, 53.34893,
    54.87195, 56.89828, 60.37057, 65.80631, 75.73663, 84.33022, 82.40794,
    84.05132, 86.21972, 84.07657, 79.09477, 72.59616, 69.73164, 62.70142,
    55.48253, 59.60514, 62.94635, 67.00214, 68.6861, 70.27246, 79.65179,
    73.4622, 47.11968,
  53.74213, 56.49059, 59.57287, 62.93986, 65.77862, 71.06311, 80.67889,
    89.92128, 92.69611, 91.5631, 90.88071, 85.53871, 77.26952, 76.8716,
    77.10579, 76.97504, 76.0731, 71.09476, 65.31828, 63.33089, 59.50417,
    58.29382, 61.25405, 64.5959, 66.17792, 65.39812, 69.07309, 74.22733,
    62.04063, 41.34515,
  64.65121, 69.28869, 73.47218, 78.04352, 81.48695, 88.38937, 92.86385,
    82.34267, 74.68069, 72.49584, 67.90735, 62.92496, 59.66474, 59.52552,
    59.95422, 61.38382, 62.45731, 61.33197, 58.76008, 58.29099, 57.73417,
    58.60254, 61.2648, 63.58159, 63.31181, 64.75171, 70.52663, 69.0941,
    54.65234, 41.33323,
  71.74127, 74.37099, 76.05339, 77.18757, 78.797, 78.44432, 67.9772,
    62.78899, 62.44683, 61.22106, 60.16083, 59.77043, 61.142, 65.61681,
    67.9604, 63.87406, 64.97456, 67.29105, 66.71465, 63.38589, 62.19775,
    65.69657, 69.56597, 69.09175, 67.04802, 72.71407, 74.86695, 63.49709,
    44.0848, 42.05915,
  74.99622, 77.71378, 74.55788, 75.15733, 76.54813, 71.19577, 57.56587,
    62.33954, 63.58992, 67.14262, 70.956, 74.92117, 74.92715, 73.87622,
    72.15071, 74.03136, 75.41161, 75.2428, 73.87769, 73.16896, 74.17431,
    72.60429, 69.75301, 65.82665, 69.31134, 76.64415, 70.45654, 50.50303,
    41.40721, 41.24893,
  76.30215, 76.43613, 77.15871, 76.91402, 80.29182, 75.6395, 69.56377,
    74.50376, 78.7473, 79.43559, 73.072, 64.40167, 63.02681, 63.38188,
    63.8319, 65.08076, 66.28779, 66.50356, 66.80347, 68.5304, 72.30705,
    69.42027, 62.69284, 61.78809, 66.8009, 65.64263, 52.1243, 41.68521,
    42.09932, 41.12288,
  84.95914, 79.64336, 87.12082, 91.73802, 87.43355, 77.93327, 79.49857,
    73.31807, 67.82085, 66.33968, 61.81387, 59.29097, 61.2211, 61.51004,
    60.10997, 60.58488, 59.9795, 60.184, 60.44609, 62.4386, 66.69633,
    66.09894, 61.9206, 67.0675, 68.51776, 56.55683, 42.35286, 44.22395,
    42.60339, 41.62714,
  104.1223, 106.5003, 108.7367, 108.4148, 106.3423, 102.5572, 85.73236,
    74.02232, 79.05862, 71.08322, 67.6973, 66.30052, 70.39188, 72.10149,
    67.64939, 59.17464, 60.63198, 60.82001, 61.17579, 63.84789, 66.9147,
    66.49006, 63.87592, 60.21024, 56.91745, 50.56727, 43.7773, 45.06926,
    43.95172, 42.48781,
  106.225, 106.8722, 105.7808, 102.44, 99.52015, 97.86806, 96.80312,
    95.96696, 89.51201, 89.83944, 93.94463, 91.76021, 89.91495, 89.53552,
    83.25435, 72.15851, 69.69041, 74.41967, 76.76888, 71.74602, 66.11559,
    61.16307, 55.8409, 49.38477, 45.78339, 44.89553, 43.67823, 43.12312,
    42.97145, 42.24553,
  100.2633, 94.31821, 91.90633, 88.98667, 88.56595, 92.46725, 97.89946,
    94.74935, 89.02367, 88.35492, 85.77367, 82.00828, 82.10222, 84.36182,
    83.86128, 82.20432, 77.00666, 73.56592, 71.39096, 66.16483, 56.25422,
    53.02945, 47.43268, 44.62792, 44.43169, 44.00687, 43.22823, 42.40098,
    41.9015, 41.51143,
  84.76071, 85.2347, 85.34174, 84.13412, 82.7737, 83.43158, 84.27579,
    80.95024, 76.29485, 72.98743, 71.91209, 69.70254, 69.3311, 72.34374,
    69.94721, 68.4009, 67.39024, 62.26041, 58.91785, 54.32763, 48.38786,
    47.89384, 44.9771, 44.17769, 44.22927, 43.84765, 43.10303, 42.40759,
    41.8256, 41.42773,
  74.08781, 72.564, 71.75925, 71.25063, 70.72276, 70.11569, 70.17558,
    70.7195, 69.27232, 66.67464, 63.40622, 66.1433, 69.89598, 67.34756,
    63.14154, 60.76092, 58.3813, 56.12383, 55.2053, 52.72113, 47.53643,
    47.7188, 45.42701, 44.27776, 44.12091, 43.99229, 42.8798, 41.92777,
    41.6128, 41.3758,
  63.54884, 63.71377, 62.95009, 63.55864, 64.01471, 64.87231, 65.66132,
    66.72336, 67.12232, 66.05762, 68.41983, 71.11947, 70.19663, 68.67244,
    64.45301, 60.47182, 56.4435, 55.62992, 56.38707, 53.37698, 47.66867,
    47.29303, 45.63336, 44.80262, 43.82715, 43.27447, 42.61588, 41.51777,
    41.36437, 41.21787,
  70.58861, 67.16673, 61.06853, 58.10158, 59.46036, 59.47702, 60.06926,
    60.70946, 60.51367, 61.81145, 64.43228, 63.24413, 58.97523, 59.37853,
    58.70363, 60.04884, 64.35822, 68.21767, 67.61285, 62.12724, 53.85666,
    48.96395, 46.25401, 45.20758, 43.82319, 43.02502, 42.43285, 41.58279,
    41.29523, 41.19231,
  70.22161, 65.47159, 58.80848, 54.95488, 55.9366, 56.06144, 56.60661,
    57.24799, 58.58856, 61.46245, 62.09108, 58.59364, 58.59599, 58.19333,
    57.76563, 58.7498, 61.71403, 65.12126, 64.99326, 62.24388, 57.18177,
    51.56873, 47.5339, 46.29179, 45.00385, 43.48245, 42.64901, 41.73038,
    41.2685, 41.21086,
  67.49857, 63.54631, 56.87413, 53.50802, 54.27181, 54.72857, 55.62459,
    56.73245, 58.36641, 60.03926, 58.66865, 56.62563, 58.68892, 58.29753,
    57.0767, 56.39376, 56.59667, 56.85313, 56.61981, 55.00523, 53.71763,
    52.82806, 50.40424, 48.19967, 46.25015, 44.159, 42.66133, 41.76983,
    41.28617, 41.21741,
  65.73694, 62.76119, 56.74059, 54.08871, 54.78797, 54.48311, 55.53509,
    56.31781, 58.11698, 58.25079, 54.93884, 53.34351, 54.35431, 53.92893,
    53.07313, 52.6909, 52.19136, 52.07515, 52.36852, 52.37066, 52.26894,
    52.00174, 51.80426, 50.48989, 47.81794, 44.58252, 42.85261, 42.02827,
    41.34971, 41.21088,
  64.29429, 62.89072, 56.45734, 54.37687, 56.23746, 56.45306, 55.6786,
    54.29953, 54.40528, 53.04259, 49.85084, 50.04287, 50.59676, 50.90712,
    50.6216, 51.12766, 51.40699, 50.82895, 50.72354, 50.68956, 50.51812,
    50.0588, 49.44424, 49.24141, 48.93922, 46.0276, 43.65966, 42.96957,
    41.99442, 41.2747,
  66.87952, 66.31862, 61.63853, 60.04184, 60.33457, 59.11273, 58.85056,
    58.13188, 59.13527, 56.91904, 54.13602, 55.78821, 57.10525, 57.76114,
    57.02219, 56.59185, 56.23104, 54.83265, 52.718, 51.46568, 50.62798,
    50.06372, 49.15824, 48.46179, 48.84234, 48.82249, 46.72078, 43.99886,
    42.96258, 41.77573,
  69.65897, 66.56052, 60.71948, 58.48247, 58.61211, 57.92365, 58.52264,
    61.06194, 64.41491, 61.75291, 58.21524, 60.20505, 61.7846, 62.47065,
    61.63699, 61.31037, 60.29871, 58.81088, 56.48415, 54.52434, 53.39915,
    52.10326, 50.09681, 48.77569, 49.24238, 50.43653, 50.20829, 46.58678,
    44.40691, 42.79892,
  71.79726, 69.49647, 64.37006, 60.49088, 59.61717, 59.28094, 61.99793,
    65.76346, 66.21443, 62.55234, 61.80759, 63.02209, 64.3743, 63.84732,
    62.21403, 61.98356, 61.47364, 60.23334, 58.23819, 56.32718, 55.28833,
    53.89727, 51.1933, 49.67609, 49.99091, 50.40549, 50.83154, 47.85594,
    43.93458, 42.5025,
  72.84573, 70.01385, 65.20572, 61.98568, 60.84276, 59.8515, 62.85658,
    64.81648, 63.98242, 62.18303, 62.89464, 63.61409, 64.22024, 63.52901,
    62.44888, 62.06174, 61.42012, 60.42537, 58.8896, 57.81068, 58.12671,
    58.41143, 56.8179, 54.6319, 53.83036, 53.74886, 53.96786, 50.79295,
    44.39818, 41.62349,
  72.91808, 70.70076, 67.72923, 66.75519, 67.16214, 66.07225, 65.95729,
    64.84872, 62.57724, 62.57917, 63.12764, 64.09389, 65.12654, 65.36897,
    65.40154, 64.98602, 63.90724, 63.11189, 62.58513, 62.42609, 61.45634,
    59.43665, 56.86708, 55.18215, 54.88115, 54.67151, 54.05215, 53.39929,
    49.58551, 43.03147,
  65.52286, 65.37483, 65.94648, 66.71528, 68.50766, 70.0224, 67.22293,
    61.85632, 60.09453, 60.35159, 60.00243, 60.47415, 61.50574, 62.76954,
    63.83953, 63.87581, 62.75175, 61.35232, 59.15887, 56.8987, 55.39849,
    54.06827, 52.41779, 51.10987, 51.03618, 50.65818, 49.54107, 48.0305,
    47.00719, 44.19999,
  61.51168, 62.07047, 62.32223, 62.08142, 64.2037, 68.1407, 68.12123,
    61.83324, 59.01506, 60.26013, 60.91775, 61.53196, 61.38431, 60.40758,
    59.15491, 57.68479, 54.74989, 52.16921, 51.10584, 49.71219, 48.36177,
    48.17504, 48.074, 47.64189, 47.25583, 46.91868, 46.06398, 44.59432,
    43.19167, 41.58879,
  41.55398, 41.47931, 41.47918, 41.4702, 41.48672, 41.53331, 41.61229,
    41.78234, 42.04208, 42.37953, 42.98866, 42.89206, 41.81021, 42.07122,
    42.18769, 41.87106, 41.8398, 41.95014, 42.1551, 42.60492, 42.75163,
    42.19167, 42.3032, 43.28916, 44.54743, 44.96903, 46.22138, 47.72208,
    43.93097, 42.30466,
  42.18206, 42.16615, 41.90298, 42.16293, 42.02465, 41.93542, 42.17927,
    42.48905, 42.88039, 43.27251, 43.63799, 43.91907, 43.95787, 43.3695,
    42.89922, 42.93608, 42.33206, 42.4768, 42.84068, 43.02544, 42.64501,
    42.71855, 44.61367, 49.27041, 53.95028, 51.29219, 46.25954, 48.96716,
    44.61772, 42.81993,
  42.22171, 42.15179, 42.14258, 42.10785, 42.00194, 42.05712, 42.20192,
    42.42757, 42.64363, 42.82038, 43.05582, 43.42611, 43.7558, 44.02945,
    43.97977, 43.09542, 43.16053, 43.91906, 44.85849, 47.12259, 51.87809,
    58.81722, 63.09587, 63.53566, 62.63115, 57.61047, 53.11327, 48.55182,
    44.63134, 43.37042,
  42.18842, 42.22195, 42.60299, 43.03589, 43.39917, 43.92337, 44.10826,
    44.18151, 44.54106, 45.0645, 45.3912, 45.79684, 45.79053, 45.42967,
    46.55539, 47.54119, 47.67128, 48.74235, 52.8934, 59.04963, 67.32193,
    69.83532, 65.0399, 64.77198, 61.12729, 59.45256, 57.91315, 50.28711,
    43.72349, 42.30682,
  43.17113, 43.24554, 44.18428, 45.00582, 45.62681, 46.00341, 46.1668,
    45.94137, 45.78365, 45.14631, 43.96181, 43.65956, 43.9496, 45.26929,
    47.40261, 50.37769, 52.78999, 55.30551, 60.93502, 67.58038, 68.48348,
    60.24721, 56.13299, 58.41509, 59.35986, 59.16896, 58.72847, 63.58181,
    62.14653, 49.30556,
  44.43844, 45.2478, 46.16445, 46.68622, 45.61946, 44.15048, 43.67206,
    43.13444, 43.62157, 45.84706, 50.35004, 60.1436, 70.01682, 70.77322,
    74.60513, 78.2806, 78.16483, 76.38445, 72.66916, 69.59518, 61.17867,
    52.01428, 55.19788, 58.02682, 61.53793, 63.2272, 65.2241, 75.26181,
    72.06895, 47.85968,
  44.68233, 45.16935, 45.87466, 46.66248, 47.30618, 50.34659, 58.74715,
    69.34641, 74.73286, 77.25362, 80.99048, 80.18173, 75.48905, 77.04481,
    78.40904, 78.52351, 77.60489, 71.67316, 64.58408, 60.83554, 55.95065,
    54.63665, 58.39697, 62.10567, 64.3844, 64.59143, 68.83525, 74.67198,
    62.7936, 41.58851,
  46.08492, 48.62261, 52.35984, 57.38754, 63.38036, 74.68736, 84.94247,
    79.68837, 75.6424, 76.13031, 73.60954, 69.17522, 65.64984, 64.84248,
    63.74441, 63.32346, 62.42254, 59.52948, 56.37886, 55.94812, 55.96323,
    57.50652, 60.53109, 63.20737, 63.47178, 65.22066, 71.09837, 70.05847,
    54.87868, 41.48233,
  55.41692, 60.77075, 65.8987, 71.29321, 78.11206, 82.21294, 74.5267,
    68.8734, 67.84983, 65.57774, 62.91068, 61.14098, 60.96458, 63.05197,
    63.63148, 59.54927, 59.88585, 61.69266, 61.81329, 59.80787, 59.26233,
    62.50641, 66.22185, 66.45608, 65.61206, 71.83745, 75.38445, 64.49232,
    44.33845, 42.04665,
  69.5401, 75.82703, 75.46981, 78.11627, 80.91442, 75.42567, 59.47789,
    61.80372, 61.42432, 62.9833, 65.56548, 68.33672, 68.09158, 67.11369,
    65.5087, 66.73677, 68.42976, 69.02223, 68.40729, 68.246, 69.37144,
    69.07609, 67.5718, 64.82173, 68.55804, 76.64651, 71.88469, 51.1656,
    41.63408, 41.60758,
  75.76785, 78.33974, 77.66883, 75.68037, 77.09052, 69.14838, 61.55122,
    67.09913, 71.54829, 74.01121, 69.52763, 62.0047, 60.59043, 60.75271,
    61.08729, 62.79713, 64.21555, 64.77599, 65.58737, 67.75072, 71.41615,
    69.45023, 64.06091, 63.78018, 69.56191, 68.89282, 54.02639, 41.95213,
    42.22961, 41.43555,
  77.92486, 69.93356, 73.7338, 77.8486, 75.77682, 69.66444, 74.84767,
    71.24521, 66.31189, 66.23361, 60.98032, 57.40756, 59.44472, 60.04764,
    59.01538, 60.24883, 60.23937, 60.78154, 61.33376, 63.26235, 67.27682,
    66.93527, 63.73841, 68.88958, 70.84782, 58.4427, 42.5943, 43.78322,
    42.61317, 41.79976,
  91.55534, 94.04176, 98.02489, 100.1112, 100.2539, 98.09219, 82.49445,
    68.93848, 73.79913, 67.1235, 63.28941, 63.27514, 67.94949, 69.88213,
    65.93846, 57.92294, 59.36596, 59.99376, 60.65426, 63.30183, 67.31177,
    68.69122, 67.00053, 62.93256, 58.54014, 50.86394, 43.32385, 44.97469,
    43.69954, 42.53938,
  98.0244, 102.2653, 103.4222, 100.7794, 97.48923, 93.89688, 90.97639,
    90.00488, 81.04271, 82.286, 88.14654, 85.92174, 84.42789, 84.38589,
    78.26009, 67.63211, 66.63377, 72.686, 76.44965, 72.64545, 68.80338,
    64.6176, 58.28454, 51.08004, 46.65021, 45.15676, 43.90763, 43.46982,
    43.11019, 42.42967,
  99.85862, 99.65558, 96.44334, 90.29564, 84.84328, 86.2205, 91.98582,
    91.95059, 86.99866, 88.06201, 85.54414, 80.17639, 79.63322, 82.08144,
    82.52255, 82.31453, 78.51205, 76.90626, 74.66375, 68.56984, 58.58086,
    54.40369, 48.17448, 44.65561, 44.51874, 44.21796, 43.49902, 42.65717,
    42.19064, 41.79092,
  92.5995, 88.19288, 85.54794, 83.40453, 83.06508, 85.35023, 86.96, 83.69626,
    79.16792, 75.06489, 73.04902, 70.99467, 71.90125, 75.9661, 74.7444,
    73.10634, 71.52022, 65.51907, 60.80781, 55.08461, 49.07401, 47.59064,
    44.55285, 43.85783, 44.26241, 44.0254, 43.23662, 42.55508, 42.01709,
    41.68598,
  81.45277, 79.44293, 79.09569, 78.70981, 77.75164, 75.81297, 74.36646,
    73.78542, 71.3937, 68.68091, 66.37543, 68.92198, 72.49158, 70.54319,
    66.02781, 62.79375, 59.53912, 56.26003, 54.22144, 51.45481, 47.00465,
    46.86239, 44.8095, 43.91566, 44.021, 44.04346, 43.05341, 42.15664,
    41.84984, 41.66784,
  73.18079, 73.25907, 71.87074, 70.83327, 69.3148, 68.63643, 68.61086,
    69.37589, 69.51785, 68.41096, 70.20366, 72.34138, 71.10535, 68.49532,
    63.47372, 59.08593, 54.78643, 53.30832, 53.52882, 51.133, 46.76825,
    46.63839, 45.11863, 44.3219, 43.77955, 43.45681, 42.78326, 41.8326,
    41.67404, 41.54768,
  77.79742, 74.2367, 67.66273, 63.86273, 64.5775, 64.58485, 65.22899,
    65.77472, 65.28047, 65.63232, 67.04245, 64.72626, 59.34653, 57.76634,
    55.33587, 55.10909, 58.22249, 61.89975, 62.21851, 58.55432, 52.29987,
    48.30465, 45.82622, 44.97367, 43.91989, 43.29185, 42.68511, 41.85272,
    41.59676, 41.52376,
  76.61696, 71.30269, 64.39059, 60.45692, 61.35966, 61.12223, 60.96539,
    60.64287, 60.48979, 61.51429, 60.62786, 56.22451, 54.87944, 53.89867,
    53.25794, 54.58428, 58.31221, 62.66772, 63.32636, 60.72736, 55.76617,
    50.54797, 47.05611, 46.06595, 44.91093, 43.69495, 42.91419, 42.00764,
    41.56241, 41.52596,
  72.40986, 68.02429, 61.21241, 57.39458, 57.457, 56.76791, 56.25484,
    56.05038, 56.53598, 57.34112, 55.74801, 53.87951, 56.09668, 56.46753,
    56.32099, 56.75546, 57.75148, 58.18276, 57.36996, 54.81192, 52.62141,
    51.28571, 49.22237, 47.57537, 45.92389, 44.22799, 42.94372, 42.04158,
    41.59118, 41.53415,
  69.03816, 65.45633, 58.74955, 55.13556, 55.06887, 54.04663, 54.3856,
    54.99661, 56.72585, 57.40902, 55.45654, 54.9287, 56.60452, 56.61874,
    55.86973, 55.15097, 53.95156, 52.89638, 52.19232, 51.40754, 50.9451,
    50.60402, 50.51348, 49.31215, 47.14124, 44.51464, 43.03902, 42.23801,
    41.66022, 41.5513,
  66.39861, 63.9428, 57.11734, 54.35687, 55.83961, 56.1337, 56.05258,
    55.67243, 56.5297, 55.90296, 53.48864, 53.57181, 53.7608, 53.25327,
    52.13982, 51.68843, 51.14568, 50.2478, 49.99268, 49.92487, 49.81398,
    49.51118, 48.92204, 48.28008, 47.81115, 45.36294, 43.41111, 42.89394,
    42.14591, 41.58705,
  67.20527, 66.18604, 61.37524, 59.59797, 60.10625, 59.2354, 59.24456,
    58.98093, 60.01108, 58.06205, 55.44921, 56.33739, 57.02726, 56.83105,
    55.66531, 55.08775, 54.57037, 53.37296, 51.74808, 50.70719, 50.08909,
    49.65327, 48.57108, 47.67424, 47.89276, 47.57128, 45.69963, 43.66416,
    42.94262, 42.00477,
  69.97154, 67.34341, 61.52122, 58.96746, 58.7678, 57.8879, 58.383, 60.41988,
    63.1785, 60.64504, 57.51073, 58.9995, 60.15573, 60.57794, 59.63681,
    59.21722, 58.50229, 57.19468, 54.99799, 53.35987, 52.51468, 51.38629,
    49.42645, 48.13416, 48.67892, 49.36702, 48.51072, 45.66127, 44.10169,
    42.84133,
  70.66462, 68.44534, 62.80597, 59.04656, 58.19302, 57.67525, 59.89404,
    63.52622, 64.32236, 61.05917, 60.51873, 61.78336, 63.09993, 62.79518,
    61.24977, 60.80333, 60.32743, 59.0577, 57.07924, 55.41025, 54.38836,
    52.85511, 50.28893, 49.09866, 49.63812, 49.54757, 49.25332, 46.86446,
    43.87915, 42.61138,
  70.75999, 68.12119, 63.01113, 59.66148, 59.03246, 58.26999, 60.89501,
    63.20272, 63.05627, 61.38631, 62.16749, 62.96461, 63.62902, 62.99799,
    61.54205, 60.84864, 60.36011, 59.30294, 57.7058, 56.60527, 56.23089,
    55.82339, 54.44027, 52.97694, 52.63318, 52.12479, 51.64957, 48.99939,
    44.00301, 41.86751,
  70.55272, 68.27909, 64.60358, 63.35492, 64.19077, 63.78878, 64.17653,
    63.74672, 62.08834, 61.96458, 62.46948, 63.22069, 64.16931, 64.19539,
    63.34412, 62.65877, 62.01537, 61.43052, 61.18103, 60.99891, 59.76747,
    57.69449, 55.24817, 53.93666, 53.72633, 53.17595, 52.1808, 51.29042,
    47.89603, 42.88779,
  64.14139, 63.93281, 64.05005, 64.46914, 66.41441, 68.17754, 66.01766,
    61.54724, 60.01031, 60.2153, 59.947, 60.27435, 61.3326, 62.45763,
    63.0328, 63.03196, 62.4766, 61.57197, 59.90416, 58.04691, 56.38938,
    54.77684, 52.95101, 51.62966, 51.43026, 50.91448, 49.74992, 48.07029,
    46.56801, 43.90703,
  60.4479, 60.91127, 61.20337, 61.15063, 63.07002, 66.50594, 66.4959,
    61.28289, 58.89346, 59.85071, 60.45303, 61.11964, 61.30773, 60.775,
    59.75875, 58.64818, 56.36363, 54.21566, 53.04694, 51.46151, 50.08903,
    49.61792, 49.2344, 48.70091, 48.12129, 47.60351, 46.50058, 44.86335,
    43.48697, 42.00512 ;

 receptor = 1, 2, 3, 4, 5, 6, 7, 8, 9 ;

 no2_conc_recp_ctl =
  31.63985, 14.40264, 31.81454, 18.16138, 13.95671, 7.219785, 25.44047,
    64.45132, 18.73225,
  67.34953, 42.34248, 68.09168, 58.15782, 48.36039, 30.06777, 64.36369,
    64.18037, 66.66003,
  65.0574, 65.00662, 66.93155, 65.22459, 65.37211, 64.98389, 66.05421,
    62.78352, 68.5452,
  61.73008, 64.09682, 64.19823, 63.83847, 62.70108, 62.02969, 64.49474,
    59.28767, 59.81551,
  59.47805, 60.71476, 60.78777, 60.42198, 57.74674, 55.70721, 62.95584,
    59.33668, 54.3748,
  61.613, 62.38839, 62.2351, 61.97882, 60.81487, 61.2836, 66.05243, 62.60542,
    59.28628,
  64.28251, 64.41595, 64.8251, 65.05736, 64.73605, 62.87738, 69.62439,
    67.69321, 64.53751,
  67.75669, 67.89587, 67.23502, 71.08678, 70.78923, 69.45512, 69.08403,
    69.39051, 67.55672,
  58.31727, 69.83437, 55.51167, 69.46463, 57.87745, 69.265, 61.80235,
    52.56347, 50.1212,
  46.87401, 66.29102, 45.73977, 60.74361, 45.6404, 60.61685, 49.69271,
    44.02885, 39.08851,
  36.73042, 54.22313, 36.08897, 52.14608, 36.63609, 47.70678, 39.37819,
    34.5997, 30.87102,
  27.63158, 48.23885, 26.53845, 41.1531, 24.57619, 38.04622, 29.51443,
    25.48495, 22.71895,
  21.29666, 37.19534, 20.11599, 33.92031, 14.76172, 27.08603, 23.2596,
    19.04246, 17.12848,
  20.6402, 38.26841, 19.52879, 29.62388, 13.45229, 20.67454, 22.31903,
    18.30339, 16.37745,
  21.01816, 39.78519, 19.78248, 29.59036, 13.2337, 19.77708, 22.6266,
    18.51625, 16.27901,
  23.96747, 51.15915, 22.36533, 31.54761, 15.36172, 21.00576, 24.58694,
    21.02692, 17.27275,
  30.55014, 78.7473, 28.21576, 41.23067, 19.67479, 29.25567, 30.05909,
    26.18474, 20.19209,
  46.24937, 71.62376, 47.08752, 64.89626, 24.791, 61.61988, 52.17236,
    36.8969, 39.80725,
  114.0698, 106.0853, 100.9665, 111.4661, 48.81997, 85.22855, 119.4085,
    89.59888, 69.856,
  91.74116, 114.075, 75.74072, 83.34864, 82.34708, 86.78671, 100.2586,
    76.81769, 62.77241,
  78.43913, 78.6936, 67.36191, 68.97374, 66.9287, 69.32494, 83.22315,
    66.69794, 55.75858,
  79.47311, 82.90139, 62.87467, 66.83922, 66.48158, 64.77215, 73.36704,
    68.07256, 59.04848,
  82.20432, 88.56595, 63.14154, 72.98743, 57.56587, 74.08781, 70.19663,
    69.75301, 58.59599,
  82.31453, 84.84328, 66.02781, 75.06489, 59.47789, 81.45277, 71.10535,
    67.5718, 54.87944 ;

 realisation = 1, 2, 3, 4, 5, 6, 7 ;

 no2_conc_grid_ens =
  7.138876, 5.89495, 6.383078, 6.462421, 6.542392, 6.653007, 6.877701,
    7.182745, 7.704432, 8.774975, 10.85496, 13.49551, 15.77814, 20.11687,
    25.1085, 30.96543, 37.708, 45.32723, 52.32591, 59.85309, 67.45981,
    73.81892, 78.35169, 81.21967, 81.87536, 79.43163, 77.78014, 80.58927,
    74.62327, 71.89901,
  5.192617, 4.210949, 4.599854, 5.153557, 5.410448, 5.585659, 5.968771,
    6.223853, 6.529876, 7.24773, 8.941141, 11.96109, 15.97234, 19.66249,
    24.44825, 31.23532, 38.76537, 45.68832, 53.06882, 61.2725, 68.55077,
    74.95367, 79.63654, 82.53423, 83.62981, 82.93416, 77.17081, 78.90222,
    74.72388, 72.5216,
  8.271354, 7.830337, 8.933871, 9.524315, 10.37959, 11.34939, 12.17687,
    12.92349, 13.4546, 13.83088, 14.56528, 16.19629, 18.88026, 22.5792,
    27.0134, 31.67291, 38.82481, 47.01468, 54.88475, 63.34074, 71.25695,
    77.66586, 82.16651, 84.35005, 84.63935, 83.96172, 83.41203, 80.36031,
    73.63993, 72.41864,
  11.02888, 11.10953, 12.73835, 13.80424, 14.41516, 14.56767, 14.70585,
    14.83484, 15.20003, 16.02045, 17.54021, 19.58351, 22.27651, 25.96145,
    30.39877, 35.28698, 41.08014, 47.31936, 54.96249, 63.46356, 71.65077,
    78.16222, 82.16693, 84.64965, 85.04211, 84.97524, 84.86726, 83.83603,
    82.32634, 73.23989,
  13.73118, 14.15354, 14.90695, 14.82667, 14.89551, 14.88385, 14.95154,
    15.02989, 15.46713, 16.54152, 18.34694, 20.91627, 23.91686, 27.58385,
    31.87658, 36.80274, 42.48069, 48.97781, 56.38588, 64.88765, 72.40742,
    77.94107, 82.07279, 84.22323, 84.84422, 84.74304, 84.45646, 85.29911,
    84.8962, 82.86357,
  13.29241, 14.39834, 15.14722, 15.3196, 15.43057, 15.40376, 15.59978,
    15.76683, 15.89944, 16.56207, 18.13635, 20.6662, 24.28384, 28.22705,
    32.75413, 38.17717, 44.66142, 51.21362, 58.61835, 66.68692, 73.67432,
    78.73559, 82.56721, 84.23605, 84.55894, 84.30342, 83.76691, 84.26209,
    84.21099, 77.22495,
  13.57656, 14.00542, 15.10632, 15.30343, 15.60864, 15.85468, 16.23267,
    16.67605, 17.09246, 17.71885, 18.98833, 20.69328, 21.34619, 26.42333,
    31.69651, 37.28823, 43.56746, 51.07143, 58.49297, 67.04183, 74.18107,
    79.499, 82.92608, 84.57094, 84.71696, 84.04195, 83.79676, 83.90819,
    83.16934, 70.11515,
  16.24004, 14.79052, 15.40424, 15.47042, 15.66552, 16.12871, 16.49152,
    15.55946, 12.71794, 16.62595, 18.24548, 20.50968, 23.44632, 27.26436,
    31.95449, 37.0753, 43.53824, 51.07782, 59.12202, 67.26811, 74.55166,
    79.98769, 83.30949, 84.61261, 84.50315, 84.25214, 84.4026, 83.95272,
    82.47375, 70.50052,
  19.01478, 16.81368, 16.76691, 16.46454, 16.32146, 16.25402, 15.29419,
    14.48344, 14.95493, 15.88825, 18.68326, 21.37957, 24.38885, 28.21153,
    32.75393, 37.16041, 43.31124, 51.4239, 59.8913, 68.07732, 75.21573,
    80.6857, 83.71301, 84.46227, 84.18395, 84.54817, 84.46671, 83.40872,
    70.97676, 71.24526,
  23.96805, 21.42944, 20.20713, 19.05248, 18.51761, 17.51181, 15.71463,
    16.02633, 16.18136, 17.12888, 19.20453, 22.62207, 26.1068, 29.08171,
    32.85547, 38.17104, 44.22869, 51.37511, 59.40848, 68.03391, 75.80747,
    81.16866, 83.22491, 83.36223, 83.76022, 84.20782, 83.83937, 77.94932,
    70.36496, 70.07198,
  28.94224, 25.73994, 25.80783, 23.42617, 22.29636, 20.45575, 18.81507,
    17.84175, 17.84915, 19.00696, 20.58015, 23.42078, 26.09458, 29.77775,
    33.99121, 38.98856, 44.82967, 51.62743, 59.14692, 67.13193, 75.51987,
    80.95486, 83.03359, 83.36452, 83.82766, 83.5442, 79.39782, 70.97705,
    71.37218, 70.19302,
  29.68075, 26.83477, 29.57512, 29.70174, 28.39459, 24.69217, 21.55295,
    18.72763, 17.74441, 18.79447, 20.6511, 23.38699, 27.36205, 30.72878,
    34.52852, 40.19705, 45.49102, 52.34279, 59.85475, 67.44515, 74.73668,
    80.70972, 82.84819, 83.82144, 84.07585, 83.16426, 71.12429, 75.64227,
    72.12975, 70.93992,
  20.10275, 21.05414, 23.53191, 26.37152, 28.12036, 27.31477, 21.17668,
    16.43847, 20.12294, 19.47872, 21.64042, 23.55689, 26.73616, 30.26358,
    34.58151, 39.17631, 45.53657, 52.60115, 60.21537, 68.08752, 75.13289,
    80.20451, 82.59928, 82.12454, 81.59592, 80.10498, 72.04095, 73.69068,
    73.14587, 71.85668,
  16.32362, 14.68464, 15.05962, 15.36828, 15.92718, 16.47488, 17.15511,
    18.48149, 17.70072, 19.20484, 21.70982, 24.8011, 27.64208, 30.6516,
    35.09706, 39.88009, 44.90746, 53.05443, 61.16228, 68.84311, 74.99986,
    79.57544, 79.77484, 75.04028, 71.68719, 71.92162, 71.39989, 70.95586,
    71.08012, 71.10255,
  17.04531, 12.22018, 15.83698, 16.02793, 16.32957, 16.50138, 16.81425,
    17.00954, 17.74663, 19.69697, 22.23005, 25.26566, 28.31668, 31.85912,
    35.22645, 39.24281, 45.7425, 51.34599, 60.13961, 68.63244, 71.92741,
    76.34595, 74.78272, 72.85966, 73.34358, 72.38354, 71.64353, 71.12508,
    70.47147, 70.3184,
  11.24889, 11.83626, 13.59836, 15.4874, 16.16144, 16.70975, 17.4126,
    17.83286, 18.74419, 21.15891, 24.54487, 27.49248, 30.52461, 32.8104,
    36.28486, 40.7098, 45.33625, 51.31598, 57.36829, 64.2462, 67.23029,
    72.18042, 72.74731, 72.8903, 72.94721, 72.32122, 71.55989, 71.06499,
    70.54594, 70.36652,
  8.199514, 6.137463, 7.739039, 9.322599, 11.21899, 13.62398, 16.088,
    16.99104, 18.54848, 21.14841, 24.29467, 27.99346, 32.42412, 35.57844,
    39.11094, 42.88815, 47.22834, 53.35255, 60.30095, 65.94884, 67.75167,
    72.42993, 73.18297, 73.0028, 72.94173, 72.56679, 71.49463, 70.48734,
    70.20651, 70.25452,
  11.46099, 7.861933, 6.779451, 7.143841, 8.483315, 9.687315, 11.08258,
    12.66936, 15.27539, 18.47913, 21.94082, 26.21426, 30.48344, 36.36199,
    41.1819, 45.21089, 49.74897, 56.44556, 64.61387, 71.80458, 71.06006,
    73.09445, 73.61892, 73.60767, 72.91904, 72.37627, 71.61313, 70.38741,
    70.05265, 70.09026,
  25.24397, 16.98601, 9.748152, 4.589466, 6.67286, 6.896639, 7.955569,
    9.221308, 10.6043, 13.17049, 17.41431, 21.19725, 24.26851, 31.7681,
    39.7598, 45.46289, 51.75349, 59.79615, 68.7363, 75.91194, 79.97339,
    77.49686, 75.53468, 75.19106, 73.71355, 72.83755, 71.98218, 70.60724,
    70.02354, 70.13338,
  24.58658, 17.15258, 10.05898, 5.114771, 6.627266, 6.926388, 7.931784,
    9.193161, 11.37497, 14.76576, 17.68622, 18.55079, 22.54597, 26.5127,
    31.80851, 38.36424, 47.18425, 57.74353, 67.16164, 74.56445, 80.00226,
    80.77436, 78.0267, 76.86356, 75.14301, 73.4761, 72.27493, 70.82085,
    70.03355, 70.16484,
  26.57431, 19.59398, 12.38902, 7.471352, 8.465275, 8.386112, 9.136183,
    10.18071, 12.2354, 14.86969, 16.36608, 18.02204, 23.20159, 27.22317,
    31.64909, 37.56567, 44.99525, 53.90236, 63.13239, 70.84377, 76.77578,
    80.65508, 80.57032, 78.71229, 76.52829, 74.21906, 72.47144, 70.92216,
    69.98717, 70.14269,
  27.76588, 23.17343, 16.15538, 12.26711, 13.81857, 13.33628, 13.95176,
    14.42197, 16.24236, 17.90454, 18.31446, 20.63103, 25.20635, 29.57319,
    34.09552, 39.95676, 46.74854, 54.58034, 62.51001, 69.35265, 74.86571,
    78.4275, 80.52152, 80.48383, 78.51775, 75.17255, 72.9362, 71.44948,
    70.1937, 70.14095,
  28.67155, 24.76015, 19.26343, 16.0994, 18.90051, 20.00496, 20.7426,
    20.89388, 22.05313, 22.87246, 23.82864, 27.72589, 32.05171, 36.53198,
    40.84324, 46.34376, 52.63985, 58.84737, 65.43407, 71.16685, 75.7461,
    78.48956, 79.45405, 79.83036, 80.15437, 77.46455, 74.20661, 72.32171,
    71.01704, 70.29646,
  28.78514, 24.73149, 21.11492, 18.67142, 20.62754, 21.15855, 22.44265,
    24.13701, 26.24358, 27.97292, 29.69728, 34.95814, 40.01375, 44.6651,
    49.01721, 54.25427, 60.22696, 65.87154, 71.31445, 76.35297, 80.03386,
    81.41489, 80.88796, 80.36597, 80.82504, 80.41177, 77.75671, 73.80257,
    72.24744, 71.0924,
  28.05332, 23.42553, 19.04671, 15.83516, 17.90856, 18.94356, 20.7028,
    22.72744, 25.05757, 26.87743, 28.58359, 33.96629, 39.42322, 44.30608,
    48.54131, 53.97647, 59.908, 66.5042, 73.02729, 78.46449, 82.24767,
    83.36215, 82.07631, 80.31268, 80.57213, 80.38444, 79.36751, 75.72707,
    72.94864, 71.9113,
  30.35221, 26.02173, 22.56537, 18.91917, 19.71288, 20.34109, 22.87486,
    25.03432, 26.91951, 28.43598, 31.54652, 35.77002, 40.93406, 45.48469,
    49.33435, 54.30486, 59.80155, 66.01234, 72.59953, 78.80157, 83.33326,
    85.26691, 83.99623, 82.31119, 81.91547, 80.77188, 79.89902, 76.83745,
    72.538, 71.31355,
  41.90601, 38.27879, 34.77126, 31.47512, 32.00849, 31.34494, 33.52884,
    35.25501, 36.16259, 37.49814, 41.14825, 45.45539, 50.12343, 53.73367,
    56.54643, 59.923, 63.67097, 68.25943, 73.69004, 78.98494, 83.05049,
    85.40849, 85.48029, 84.35891, 83.72003, 82.71645, 82.23769, 79.97301,
    74.34415, 70.93777,
  60.26619, 58.70781, 55.84294, 54.37965, 55.50919, 56.00843, 55.36275,
    54.8214, 53.87102, 54.94682, 56.51288, 59.26625, 62.74636, 65.46236,
    67.11285, 68.79411, 70.03368, 72.22272, 75.66514, 79.54751, 81.39595,
    81.84238, 81.12499, 80.36655, 80.50678, 80.17111, 79.74167, 79.48942,
    77.39925, 72.50415,
  69.53883, 70.02304, 71.95985, 72.89028, 73.91319, 75.18822, 74.82116,
    70.43237, 68.91058, 69.57043, 69.42066, 69.5977, 70.278, 71.31897,
    72.12154, 72.6493, 72.68737, 72.80978, 73.4284, 74.012, 75.20426,
    76.54414, 76.77705, 76.06481, 76.32996, 76.28204, 75.62399, 74.07417,
    73.45796, 72.54285,
  74.62774, 75.147, 75.60657, 75.48273, 76.54342, 78.94859, 79.50328,
    75.91915, 73.68488, 74.60679, 75.23739, 75.71652, 75.69964, 75.41543,
    74.95987, 74.52296, 73.26183, 71.82771, 71.70296, 71.87486, 71.6504,
    72.49212, 73.34879, 73.67646, 73.65378, 74.00999, 73.59039, 72.32301,
    71.23876, 70.35967,
  32.19352, 34.84146, 38.18501, 41.90523, 45.88387, 49.85566, 53.75805,
    57.81804, 62.17168, 66.64893, 71.1581, 75.0986, 78.04939, 80.42569,
    82.01114, 82.85065, 83.19006, 83.31479, 83.28615, 83.14663, 82.66016,
    81.7331, 80.78153, 80.01382, 79.23248, 78.07845, 69.12779, 72.18422,
    68.0634, 65.16984,
  31.12523, 33.82272, 37.33268, 41.22507, 45.53577, 50.16961, 54.76567,
    59.04859, 63.252, 67.68948, 72.16557, 76.30457, 79.58644, 81.68164,
    82.8914, 83.46217, 83.5377, 83.56897, 83.59473, 83.65148, 83.52768,
    83.18845, 82.47114, 81.73416, 81.1272, 79.58685, 76.54243, 70.76063,
    67.4575, 65.49843,
  32.51788, 35.07827, 38.42842, 42.07816, 45.86591, 50.15176, 55.17138,
    60.04744, 64.5509, 68.87117, 72.91701, 76.81985, 80.10642, 82.31434,
    83.51078, 83.77018, 83.62926, 83.51607, 83.45622, 83.28876, 83.40787,
    83.49529, 83.05157, 82.33839, 81.4464, 80.72233, 79.89641, 78.23035,
    68.07373, 65.0954,
  33.31326, 36.13189, 40.12491, 43.47976, 46.76994, 50.37026, 54.70456,
    59.72313, 64.78513, 69.58115, 73.72755, 77.39089, 80.68376, 82.90524,
    84.06308, 84.46275, 84.19623, 83.75925, 83.75253, 83.62389, 83.51304,
    82.84305, 81.6333, 81.47339, 80.71786, 80.71923, 80.91341, 80.13303,
    78.3813, 68.29421,
  34.05757, 37.09662, 41.04627, 45.12753, 48.58683, 51.82506, 55.11525,
    59.66385, 64.28466, 69.29073, 73.77332, 77.53585, 81.05267, 83.53515,
    84.85184, 85.26382, 84.95332, 84.36181, 84.06968, 83.90534, 83.23514,
    81.79553, 81.1441, 80.85994, 80.5393, 80.12078, 80.02257, 81.06782,
    80.66704, 78.20505,
  35.0979, 37.9147, 41.72269, 45.85547, 50.013, 53.44644, 56.40033, 60.77195,
    64.78398, 68.94884, 73.21719, 77.16706, 80.95184, 83.488, 85.1468,
    85.8661, 85.51624, 84.87226, 84.17286, 83.73079, 82.89439, 81.48637,
    81.32691, 80.93704, 80.47916, 80.02678, 79.55367, 80.05857, 79.88596,
    70.4443,
  38.18232, 39.73389, 42.82714, 46.32267, 50.31563, 54.11847, 57.51672,
    61.76762, 66.06673, 69.92636, 73.76151, 76.86233, 78.95432, 81.58416,
    83.33421, 84.32022, 84.67743, 84.11338, 82.99569, 82.59399, 82.15765,
    81.60796, 81.2413, 81.04059, 80.60973, 80.04104, 79.82179, 79.78516,
    78.8229, 63.42558,
  43.85385, 44.28988, 45.92794, 48.13651, 51.24189, 55.31606, 59.06306,
    61.51814, 64.86433, 68.81857, 72.37885, 75.68977, 78.69706, 81.34226,
    83.14884, 84.06974, 84.64883, 84.65005, 83.91678, 82.96431, 82.18096,
    81.54281, 81.09864, 80.72386, 80.07936, 80.00165, 80.02509, 79.38298,
    77.77184, 63.86363,
  50.21322, 51.42972, 52.05237, 52.82598, 54.42482, 57.10663, 59.14582,
    62.32317, 66.31173, 69.99767, 73.29296, 76.25979, 78.69736, 81.04134,
    82.97573, 83.60921, 84.19976, 84.82214, 84.95073, 83.99571, 82.84639,
    81.78439, 80.85732, 80.04304, 79.45889, 79.89751, 79.91393, 78.76133,
    63.6861, 64.62683,
  53.69316, 57.43819, 59.22548, 59.67643, 59.79401, 60.2882, 61.01787,
    63.84664, 67.26743, 71.11657, 74.17574, 77.04129, 79.09632, 80.53461,
    81.61098, 82.74469, 83.3327, 83.68481, 84.00107, 83.8456, 83.49583,
    82.12049, 80.52858, 79.24622, 79.12514, 79.25141, 78.86149, 71.52469,
    63.88684, 63.50738,
  52.62323, 56.67737, 62.08529, 64.7752, 65.71368, 65.32003, 65.50632,
    66.73396, 68.67395, 72.61279, 75.28668, 77.30418, 79.05206, 80.36559,
    81.30106, 82.01508, 82.42976, 82.65843, 82.83482, 82.78976, 83.17419,
    82.15122, 80.27417, 79.57282, 79.61631, 78.93959, 74.30801, 65.35274,
    65.09474, 63.81974,
  48.76488, 49.76059, 58.3843, 65.06065, 70.56107, 70.35117, 68.7541,
    67.68966, 70.20038, 72.85414, 75.86701, 78.07494, 80.51932, 81.72912,
    82.08762, 82.27009, 82.74578, 82.91818, 82.81838, 82.45749, 82.77724,
    82.19069, 80.2086, 79.47517, 79.3791, 78.50799, 63.94902, 70.04381,
    66.08341, 64.67056,
  42.09577, 45.53299, 49.77451, 56.96427, 64.78746, 70.36735, 69.14665,
    66.54628, 73.18054, 74.70295, 77.87575, 79.85435, 82.14005, 83.65058,
    83.88525, 82.61482, 82.99899, 83.37042, 83.31046, 82.60359, 82.4811,
    81.93179, 80.40945, 75.51174, 73.12941, 74.30916, 64.86701, 66.29986,
    66.67203, 65.55905,
  40.25054, 42.73668, 45.51621, 49.49569, 53.86996, 58.27855, 63.63778,
    69.54202, 71.82708, 75.35994, 78.94397, 81.87291, 83.58311, 84.97359,
    85.15567, 84.08849, 83.29324, 83.5903, 83.82298, 82.67406, 81.5602,
    80.63766, 77.41785, 70.12249, 64.82346, 64.7425, 64.88401, 64.05633,
    64.1005, 64.44147,
  38.42778, 36.54152, 44.63875, 48.90455, 52.97182, 57.6548, 61.6756,
    65.94302, 71.23476, 75.44915, 78.75361, 81.42625, 83.66271, 85.48376,
    85.94078, 85.94411, 84.71558, 83.55784, 82.94539, 82.26721, 76.49698,
    76.16066, 71.23174, 67.19495, 67.28705, 65.58177, 64.87048, 64.43372,
    63.80133, 63.71749,
  32.92313, 35.91483, 39.61174, 44.49715, 49.96665, 55.06772, 59.64688,
    63.91106, 68.84962, 74.09569, 78.13239, 81.09315, 83.68893, 85.84793,
    86.81008, 86.78343, 86.42927, 84.99299, 82.79285, 78.47313, 74.21402,
    72.94907, 69.66067, 67.5396, 66.66159, 65.45899, 64.56071, 64.14003,
    63.85977, 63.778,
  36.84403, 36.01102, 39.87817, 43.63947, 48.0293, 52.99195, 58.17505,
    63.19091, 67.23126, 71.99416, 76.31316, 80.00378, 83.52053, 85.4591,
    86.70657, 87.7695, 88.22414, 87.778, 86.20789, 83.80103, 75.99819,
    73.85319, 70.77481, 68.22141, 66.96503, 65.89236, 64.6357, 63.7959,
    63.65788, 63.70064,
  47.81506, 43.465, 42.90787, 45.21368, 50.12992, 54.34512, 58.83081,
    63.4739, 67.72041, 71.51224, 75.99009, 79.68858, 82.19931, 84.10587,
    85.13443, 86.56173, 88.27673, 89.2734, 89.03455, 87.01017, 82.68166,
    75.51495, 71.74102, 69.55399, 67.37436, 66.28429, 65.09442, 63.84953,
    63.56455, 63.58684,
  57.75742, 54.71705, 50.60791, 46.3367, 52.04082, 55.44313, 60.47942,
    64.77661, 69.62524, 73.84826, 78.14086, 80.4184, 80.12305, 80.48909,
    81.34003, 83.51668, 86.38995, 88.0304, 88.72494, 88.3558, 86.33936,
    80.82991, 73.60201, 71.65516, 68.7651, 67.2055, 65.87722, 64.15715,
    63.58765, 63.63223,
  56.96697, 55.25614, 52.7566, 50.26519, 55.31347, 58.71245, 63.0102,
    67.89513, 72.76234, 77.22374, 80.45176, 82.69382, 84.78162, 84.66177,
    82.97875, 81.84299, 82.5459, 84.7038, 85.70111, 85.66224, 85.02579,
    82.93943, 76.42754, 73.18055, 70.61653, 68.16872, 66.47195, 64.46713,
    63.52777, 63.67185,
  59.18129, 57.03708, 54.60363, 54.26047, 58.84566, 62.32956, 66.97655,
    71.25479, 75.52471, 79.57187, 82.69514, 84.16552, 87.0739, 88.23019,
    87.36879, 86.59867, 85.70921, 85.44141, 84.77939, 82.79688, 81.79922,
    81.0137, 78.43546, 74.95479, 72.15678, 69.19329, 66.90792, 64.75175,
    63.52402, 63.612,
  64.69028, 62.21358, 59.38868, 58.78456, 63.21331, 66.39867, 70.3936,
    74.45563, 78.71773, 82.78934, 86.12541, 88.61196, 90.46015, 91.45654,
    91.57548, 90.99724, 89.5015, 88.11912, 86.83723, 84.54374, 81.79193,
    79.56889, 78.46415, 76.45309, 74.19933, 70.44144, 67.50188, 65.68248,
    63.94573, 63.6442,
  74.52516, 71.76389, 67.98411, 66.6928, 70.27302, 73.06932, 76.47639,
    79.92296, 83.50111, 86.87945, 90.14848, 93.28581, 95.53391, 96.2562,
    95.96394, 95.36823, 94.43154, 93.07587, 91.01053, 88.05528, 85.26531,
    81.66261, 78.8461, 76.69673, 75.87863, 72.72346, 68.91008, 66.63404,
    65.17597, 64.00598,
  85.65954, 82.42986, 78.36256, 76.42925, 78.62997, 79.87435, 82.37375,
    85.4412, 88.85643, 91.17302, 93.5406, 97.00068, 100.2527, 101.2404,
    100.52, 99.91209, 98.99548, 97.55383, 95.41623, 93.18815, 90.28692,
    86.4195, 81.47418, 78.17586, 77.40627, 75.66042, 72.31857, 67.97459,
    66.35959, 65.02232,
  93.72775, 89.81348, 84.47859, 81.10394, 82.89126, 83.37479, 84.75973,
    87.14761, 89.98779, 91.33356, 92.77346, 95.48763, 98.47984, 99.7036,
    98.61829, 98.26729, 97.59441, 96.51365, 94.88656, 93.32716, 91.08304,
    87.55897, 82.33035, 78.60553, 77.7724, 76.28701, 74.27872, 69.72328,
    66.50555, 65.56568,
  96.209, 91.57504, 86.67081, 82.00359, 82.06333, 81.34765, 83.72768,
    86.48498, 88.266, 87.56375, 89.29484, 92.31322, 95.34336, 96.34618,
    95.13606, 94.81083, 94.02314, 92.93223, 91.37267, 90.04291, 88.57066,
    86.55716, 81.89777, 78.39564, 77.84666, 76.42818, 75.25006, 71.81503,
    66.60762, 64.93633,
  93.61085, 90.24655, 85.5598, 80.35035, 80.33346, 78.25644, 79.00448,
    80.49288, 80.52098, 79.62545, 81.34454, 84.49645, 88.71759, 90.41717,
    89.2551, 88.63155, 87.56253, 86.29261, 85.49381, 84.96956, 84.34711,
    82.81158, 79.91095, 77.08218, 76.5327, 75.43117, 75.3355, 73.83075,
    68.73699, 64.99392,
  86.79823, 85.00063, 81.01269, 78.13144, 79.12921, 78.1403, 76.69141,
    75.68658, 74.32387, 73.82893, 73.8313, 75.366, 78.32204, 80.2802,
    80.2603, 80.29721, 78.99729, 77.82266, 77.58444, 78.47913, 78.39052,
    77.55611, 75.10781, 73.45557, 73.23469, 72.37415, 71.53644, 71.23179,
    70.0644, 66.15443,
  70.67422, 71.27539, 72.7834, 74.08058, 75.19592, 76.71848, 74.52193,
    71.01179, 69.56862, 70.04556, 69.67936, 69.18623, 69.09138, 69.8524,
    70.41595, 70.54482, 70.06038, 69.12981, 68.4389, 68.17909, 68.65057,
    69.87567, 70.35769, 69.57099, 69.75602, 69.46952, 68.66515, 66.84675,
    65.97359, 65.60281,
  67.87184, 68.06453, 68.63477, 68.61923, 68.98438, 70.32799, 70.74304,
    68.3455, 66.84276, 67.54365, 67.91741, 67.991, 67.59893, 67.32146,
    67.22264, 67.11718, 66.38911, 65.16601, 64.91508, 64.82864, 64.55198,
    65.10197, 66.00956, 66.557, 66.57866, 66.78046, 66.5733, 65.51225,
    64.52267, 63.776,
  74.85323, 76.99358, 78.14316, 79.39751, 80.11197, 80.50085, 80.73907,
    80.76842, 80.47814, 80.19428, 80.03432, 79.68105, 79.10403, 78.56561,
    78.2406, 78.0456, 77.92133, 77.95845, 77.98867, 77.63831, 76.82081,
    75.94428, 75.2049, 74.59673, 74.10014, 72.11267, 66.35645, 68.70972,
    65.87106, 63.81232,
  74.83154, 77.00228, 78.15006, 79.42809, 80.21001, 80.66917, 81.00678,
    81.10589, 80.8891, 80.72962, 80.57858, 80.17945, 79.56458, 79.06711,
    78.47773, 78.07634, 77.89021, 77.85789, 78.04015, 77.99557, 77.65369,
    77.20622, 76.6288, 76.19533, 75.63821, 74.2101, 70.08216, 66.82301,
    65.33852, 63.82605,
  74.98872, 77.03558, 78.13852, 79.37264, 80.19811, 80.7441, 80.9381,
    80.9127, 80.77833, 80.7171, 80.67111, 80.35918, 79.85783, 79.36536,
    78.91624, 78.377, 77.84511, 77.6378, 77.58633, 77.4959, 77.48615,
    77.48966, 77.30119, 76.92732, 76.24393, 75.35431, 74.36587, 73.03613,
    65.44214, 63.73965,
  75.17596, 77.13471, 78.23507, 79.45795, 80.35571, 81.04296, 81.21765,
    80.9882, 80.76186, 80.60465, 80.60709, 80.72095, 80.50983, 79.96163,
    79.46233, 79.03529, 78.38505, 77.85575, 77.52546, 77.29848, 77.1797,
    76.72241, 75.92582, 76.05088, 75.63189, 75.79517, 75.65681, 74.87473,
    73.69102, 66.49932,
  75.45931, 77.31658, 78.40791, 79.40266, 80.12144, 80.92786, 81.42963,
    81.30101, 80.98807, 80.57307, 80.39948, 80.81946, 81.14142, 80.79949,
    80.32264, 79.80822, 79.20287, 78.38792, 77.89701, 77.45592, 76.69359,
    75.89046, 75.47861, 75.53587, 75.46527, 75.16811, 75.28949, 76.34846,
    75.9633, 73.97007,
  76.16895, 77.70419, 78.82692, 79.69681, 80.16811, 80.84252, 81.63995,
    81.77617, 81.60175, 81.26803, 80.96584, 81.07944, 81.46527, 81.037,
    80.85605, 80.48181, 79.44561, 78.79086, 78.25258, 77.58999, 76.75135,
    75.54768, 75.66417, 75.56329, 75.28368, 74.94903, 74.7453, 75.22992,
    75.28772, 69.45558,
  78.15939, 78.65795, 79.60828, 80.40765, 80.85269, 81.25769, 81.65926,
    81.63171, 81.66222, 81.40948, 81.37854, 80.73109, 79.63503, 79.6293,
    79.29661, 79.07691, 78.86931, 77.95963, 76.99489, 76.65048, 76.12859,
    75.65813, 75.48675, 75.55744, 75.36565, 74.96353, 74.89719, 74.97338,
    74.20669, 62.47532,
  82.44243, 81.416, 81.32083, 81.64842, 81.89796, 82.22243, 82.09309,
    80.64518, 79.68347, 79.59747, 79.60069, 79.54095, 79.45454, 79.45036,
    79.40974, 79.27343, 79.05692, 78.57314, 77.82365, 77.03136, 76.29295,
    75.58799, 75.3138, 75.11445, 74.80997, 74.9799, 75.09914, 74.50715,
    73.27054, 62.79051,
  88.17149, 87.31686, 85.3383, 84.29749, 83.56332, 82.90378, 81.27157,
    81.0714, 80.68801, 79.9922, 79.59563, 79.26669, 78.93884, 78.84121,
    79.0169, 78.89098, 78.91468, 79.02538, 78.95437, 78.12537, 77.01656,
    76.02277, 75.22116, 74.48749, 74.21978, 74.71612, 74.98083, 74.0586,
    62.69365, 63.41199,
  91.46429, 93.35794, 91.85767, 89.61491, 87.3204, 84.79627, 82.1398,
    82.05164, 81.59338, 80.8978, 79.80421, 79.08147, 78.33712, 77.9538,
    77.73751, 77.78054, 77.88398, 78.10561, 78.33154, 78.28423, 77.77347,
    76.55164, 75.23991, 74.17717, 74.12589, 74.292, 74.16899, 69.13116,
    62.77941, 62.78031,
  89.41779, 92.7026, 96.04714, 95.57603, 93.36469, 88.68397, 85.35074,
    83.49265, 82.37357, 82.22985, 80.53562, 78.79696, 78.19308, 77.62903,
    77.12078, 76.97372, 76.55703, 75.37057, 75.64754, 77.22054, 77.55302,
    76.66909, 75.09039, 74.54838, 74.92889, 74.61583, 72.46523, 63.76449,
    63.88303, 62.95361,
  85.13646, 85.85455, 91.59954, 95.7345, 96.82803, 93.27069, 88.25484,
    84.49928, 83.38175, 82.68436, 81.51717, 80.28345, 79.70007, 79.08031,
    77.97967, 77.24603, 77.19243, 77.09088, 76.89771, 76.65114, 77.00479,
    76.43051, 74.93773, 74.34048, 74.5338, 74.11175, 63.08351, 68.33464,
    64.59475, 63.59936,
  79.19463, 81.47982, 83.26347, 86.79705, 90.3362, 91.93673, 87.15547,
    83.43482, 85.43414, 84.12521, 83.36695, 82.1015, 81.62709, 81.01526,
    79.64958, 77.61897, 77.61557, 77.64138, 77.34885, 76.67313, 76.63736,
    76.2794, 75.01246, 72.29732, 70.87559, 72.42768, 63.61868, 65.27377,
    65.47233, 64.37293,
  79.50813, 80.68649, 80.72219, 78.59685, 77.77178, 81.55511, 83.4944,
    84.88859, 83.1694, 83.93183, 84.16756, 83.23953, 82.52332, 82.00558,
    80.52824, 78.74951, 77.88293, 78.00435, 78.10129, 77.05138, 76.07374,
    75.25813, 72.0563, 66.48198, 62.93975, 63.51554, 63.86159, 63.2469,
    63.38457, 63.56303,
  79.76377, 78.83016, 81.75383, 81.90538, 81.96887, 82.22613, 82.675,
    82.61688, 82.38676, 82.12629, 82.20546, 82.0797, 82.17506, 81.85956,
    80.99131, 80.24696, 78.78352, 78.09132, 77.75699, 76.81714, 71.21455,
    70.96207, 67.53719, 64.21426, 64.98287, 64.40373, 63.96023, 63.56114,
    62.96157, 62.88265,
  76.48595, 78.94052, 79.87615, 80.95064, 81.22035, 82.78244, 83.05012,
    82.90846, 82.18197, 81.53499, 81.42201, 81.69505, 82.13202, 82.74355,
    82.00646, 80.96621, 80.34508, 79.20457, 74.57941, 71.83635, 69.21507,
    68.14534, 65.89674, 64.74255, 64.61765, 64.26187, 63.71084, 63.2467,
    62.94837, 62.91697,
  80.45194, 79.94428, 80.75013, 81.77097, 82.18848, 82.01443, 82.37824,
    83.62843, 83.11352, 82.0571, 81.33485, 81.53557, 82.34597, 82.53346,
    82.43535, 82.60722, 82.58453, 81.96767, 80.30141, 76.37639, 70.54136,
    69.14502, 67.13622, 65.62671, 65.2105, 64.6209, 63.68012, 62.91825,
    62.8252, 62.8807,
  88.60719, 86.06547, 83.2188, 82.97198, 83.93413, 83.84838, 83.9384,
    83.7134, 84.03802, 82.60379, 82.42502, 82.21886, 81.67593, 81.07048,
    80.90912, 81.88554, 83.18324, 83.82973, 83.27183, 81.21864, 76.24867,
    70.78077, 68.3166, 67.13368, 65.99915, 65.26371, 64.01153, 63.00347,
    62.77704, 62.84246,
  97.6357, 93.87888, 88.76888, 83.07533, 85.36915, 84.81252, 84.60544,
    84.59065, 83.6964, 83.88873, 84.04845, 82.73649, 79.44, 77.08562,
    76.37112, 78.02518, 81.14879, 82.45278, 83.00051, 82.73209, 80.75402,
    75.24158, 69.88436, 69.18359, 67.28378, 66.16965, 64.94585, 63.21672,
    62.81798, 62.84165,
  96.55251, 93.78751, 88.72631, 84.28967, 86.26376, 86.16875, 86.26437,
    85.68714, 85.62355, 85.81362, 85.96692, 85.33829, 84.88847, 81.59792,
    78.37117, 76.72208, 76.86494, 78.67868, 79.56519, 80.09777, 79.39011,
    77.12222, 72.16926, 70.27196, 68.74394, 66.97491, 65.47911, 63.586,
    62.76093, 62.91712,
  96.17904, 93.5222, 88.22125, 83.81463, 86.05889, 86.37562, 87.01282,
    87.40527, 87.8631, 87.32265, 85.97884, 84.51596, 85.08611, 84.43442,
    82.50175, 81.43427, 80.72868, 80.527, 79.76805, 77.62897, 76.36766,
    75.6925, 74.03071, 71.56039, 69.83965, 67.54028, 65.76386, 63.77763,
    62.73067, 62.80833,
  94.95273, 92.85758, 86.66465, 82.47751, 85.15639, 85.78402, 87.46427,
    88.70521, 89.93618, 90.45004, 89.41798, 87.53622, 86.90062, 86.07941,
    84.89212, 84.03172, 83.34658, 82.78534, 82.19804, 79.79036, 76.73371,
    74.74125, 74.60335, 72.3748, 71.1358, 68.56233, 66.46409, 64.50101,
    62.96607, 62.80053,
  93.41808, 90.78841, 84.69417, 80.31699, 83.47227, 84.72522, 86.86641,
    88.55613, 90.34501, 91.70819, 92.08728, 91.89469, 91.24751, 90.72694,
    89.81312, 88.9641, 88.17892, 86.86994, 85.3347, 83.21483, 80.34978,
    77.04115, 75.34901, 73.03472, 72.33717, 70.44777, 67.76705, 65.41228,
    63.99057, 63.09422,
  92.23361, 89.24201, 82.87047, 79.45807, 81.08033, 82.21341, 84.6899,
    87.28391, 90.01472, 91.53918, 92.49902, 93.70458, 94.97806, 95.3842,
    94.17595, 93.28562, 92.36022, 91.19968, 89.34769, 87.37544, 85.25504,
    82.16112, 78.007, 75.4436, 74.37267, 72.98615, 70.64766, 66.80107,
    65.12189, 63.92595,
  90.99994, 87.80734, 80.48255, 76.21573, 77.10478, 77.43642, 79.94563,
    83.77915, 87.36546, 88.30463, 89.1322, 90.92085, 93.3984, 94.52398,
    93.27556, 92.47007, 91.5703, 90.28018, 88.75183, 87.40758, 85.62714,
    82.91817, 78.98682, 76.14404, 75.43865, 73.97698, 72.22095, 68.01661,
    65.16816, 64.25184,
  89.69474, 86.29137, 81.12615, 76.07748, 75.8909, 75.11525, 77.01944,
    80.2851, 82.84879, 82.93537, 84.93543, 87.66029, 90.26395, 91.2955,
    90.30482, 89.70229, 88.86159, 87.52338, 86.51866, 85.53827, 83.96651,
    82.0624, 78.61717, 76.03102, 75.75844, 74.30637, 72.94312, 69.61522,
    65.34954, 63.88682,
  86.66882, 84.1153, 80.39802, 75.83078, 75.82435, 74.24496, 74.74577,
    76.23141, 77.25616, 77.13064, 79.04199, 82.11815, 85.2832, 86.49205,
    85.78118, 85.47913, 84.67269, 83.4715, 82.7975, 82.24203, 81.25716,
    79.65926, 77.2411, 75.17897, 74.67001, 73.68136, 73.14666, 71.3287,
    67.07327, 64.02036,
  81.26574, 80.20345, 77.31972, 74.97171, 76.02014, 75.27812, 74.03944,
    73.28876, 72.56545, 72.47044, 72.9045, 74.54302, 77.45672, 79.007,
    79.14486, 78.86222, 77.42086, 76.09174, 75.54031, 76.36221, 76.57243,
    75.82305, 73.62383, 72.01096, 72.02658, 71.18411, 70.36102, 69.70551,
    68.37743, 64.92855,
  68.7411, 69.6798, 71.0473, 71.82957, 72.74409, 74.25427, 72.70546,
    69.56303, 68.40716, 68.77575, 68.62749, 68.14203, 68.01436, 68.718,
    69.03817, 69.29681, 68.79033, 67.70963, 67.09702, 67.02363, 67.659,
    68.8513, 69.25367, 68.38513, 68.31223, 68.2672, 67.62294, 66.00884,
    65.03881, 64.612,
  66.03873, 66.42089, 67.03232, 66.88605, 67.41722, 68.76595, 69.15408,
    67.15215, 65.95593, 66.58265, 66.82996, 66.67146, 66.24837, 65.88231,
    65.88237, 65.81056, 65.23479, 64.21957, 63.94227, 63.92645, 63.6809,
    64.25961, 65.20644, 65.58155, 65.42843, 65.55649, 65.40994, 64.47979,
    63.72635, 63.0163,
  77.495, 76.97523, 76.91204, 76.78163, 76.54018, 76.3648, 76.19523,
    75.99678, 75.92307, 76.06174, 76.33639, 76.57798, 76.80607, 77.35811,
    78.12135, 79.07146, 80.18864, 81.63097, 83.27037, 84.99514, 86.48473,
    84.26709, 81.97957, 80.24979, 77.66457, 73.19107, 70.13624, 72.06314,
    69.225, 67.16193,
  77.26481, 76.77336, 76.67767, 76.47855, 76.16266, 75.91924, 75.78791,
    75.64892, 75.66192, 75.78253, 75.99619, 76.30956, 76.72965, 77.29452,
    78.03199, 79.05111, 80.11346, 81.51761, 83.26656, 85.2409, 87.13518,
    88.49097, 89.09808, 89.44067, 89.23293, 81.89379, 71.07257, 69.70146,
    68.93684, 67.31348,
  77.41547, 77.11126, 77.16246, 76.89818, 76.55448, 76.22723, 75.99379,
    75.91224, 75.96391, 76.12648, 76.42214, 76.87602, 77.37973, 77.97434,
    78.72456, 79.59505, 80.47932, 81.40762, 83.28079, 85.14545, 87.34937,
    89.23901, 90.18269, 90.39841, 89.80719, 88.53336, 87.53332, 73.37852,
    68.17916, 67.34144,
  77.15339, 76.8637, 76.98385, 76.96529, 76.797, 76.57764, 76.32782,
    76.11038, 76.09376, 76.28143, 76.76248, 77.43957, 78.05899, 78.61157,
    79.24616, 79.98023, 80.88024, 82.02036, 83.52945, 85.26358, 86.98315,
    88.39357, 85.08303, 88.91879, 89.31107, 89.29244, 88.6532, 88.11868,
    78.35823, 69.28844,
  77.14243, 76.61604, 76.6479, 76.64475, 76.66344, 76.81977, 76.97016,
    76.6852, 76.48907, 76.55299, 77.20257, 78.12994, 79.09254, 79.79725,
    80.48245, 81.15546, 81.6188, 82.11545, 83.52335, 85.42962, 86.61416,
    82.42496, 80.08717, 82.16663, 84.21201, 87.46603, 88.8207, 89.73899,
    89.80971, 79.74202,
  77.29229, 76.69376, 76.55344, 76.32, 76.16037, 76.6141, 77.46304, 77.53568,
    77.24942, 77.03799, 77.3159, 78.24416, 79.55757, 80.33859, 81.48866,
    82.6053, 82.89294, 82.87251, 83.22614, 84.73815, 86.02395, 78.9959,
    83.68372, 83.28794, 83.16973, 82.56673, 82.75397, 88.85198, 88.98077,
    73.32865,
  77.78049, 76.93587, 76.81953, 76.37487, 76.0775, 76.51101, 77.29421,
    77.53613, 77.65885, 77.62546, 77.84169, 77.71236, 77.49772, 78.60262,
    79.82005, 80.34382, 81.44713, 81.86508, 81.80406, 82.80991, 81.59465,
    80.75675, 83.58969, 86.43179, 87.43129, 86.87688, 86.95808, 88.99788,
    85.45924, 66.04928,
  79.35195, 77.71333, 77.37173, 76.8512, 76.68737, 76.88179, 76.91409,
    75.7425, 75.17548, 75.71093, 76.1619, 76.62695, 77.31594, 78.18261,
    79.1815, 80.21255, 80.97343, 81.01042, 80.28401, 79.96188, 80.10664,
    80.73646, 82.50814, 85.21803, 88.00056, 89.30109, 89.3074, 88.63033,
    79.82458, 66.2082,
  83.00654, 80.67935, 79.07467, 78.11817, 77.53778, 76.98917, 75.65961,
    75.52697, 75.63092, 75.755, 76.20988, 76.65581, 77.25124, 78.34969,
    79.49518, 80.30378, 81.58625, 83.09039, 84.36086, 85.22358, 84.47636,
    84.23299, 83.97441, 82.94068, 84.41544, 89.31293, 89.589, 87.52161,
    66.25984, 66.91769,
  87.44889, 86.16123, 83.74468, 81.5955, 80.0598, 78.09467, 76.07831,
    76.29533, 76.33261, 76.64455, 76.89215, 77.19896, 76.65608, 75.90173,
    75.92667, 77.22163, 79.0255, 80.86663, 82.88216, 85.01089, 87.19888,
    87.51989, 86.76813, 85.39035, 85.73029, 86.58627, 84.98668, 72.93343,
    66.23834, 66.33176,
  89.53708, 89.34393, 90.51984, 87.64993, 85.25703, 81.35425, 79.01756,
    77.76807, 77.37984, 78.2191, 78.03075, 77.66805, 77.8282, 76.12438,
    74.56155, 74.75597, 74.56817, 75.02234, 76.50771, 79.06953, 82.82931,
    84.38828, 84.66599, 88.55958, 89.29482, 88.95112, 74.70643, 66.69508,
    67.33709, 66.47132,
  87.93871, 87.26002, 90.74243, 92.34201, 90.73378, 86.5845, 82.34354,
    78.99473, 77.74273, 78.27162, 78.16079, 78.02736, 78.95255, 79.34385,
    79.35185, 78.58133, 78.69631, 77.44067, 76.61178, 77.2113, 80.51461,
    81.95264, 80.20131, 82.32935, 88.75339, 87.57169, 66.73672, 71.12691,
    67.86716, 66.97032,
  79.69514, 81.14162, 82.9612, 85.53636, 87.73656, 87.66759, 82.01598,
    77.70087, 79.87218, 79.01965, 79.09431, 78.88483, 79.68597, 80.2894,
    80.30558, 80.18169, 81.70691, 83.62971, 84.99483, 81.16596, 82.43267,
    84.18086, 81.57588, 75.3825, 74.11219, 74.98303, 67.12428, 68.84481,
    68.75122, 67.65177,
  79.12032, 78.17882, 77.81214, 76.64067, 76.63235, 77.60004, 79.0749,
    79.98624, 78.66206, 79.26488, 79.78313, 79.92205, 80.08555, 80.46286,
    80.52965, 80.23732, 80.78731, 83.08348, 85.30492, 86.53447, 84.12325,
    80.80502, 72.80205, 69.28516, 66.8265, 67.13223, 67.15958, 66.72658,
    66.97433, 67.00993,
  80.72731, 80.25492, 79.36026, 78.27316, 77.58305, 77.76668, 78.39929,
    78.59534, 78.75005, 79.05273, 79.33839, 79.45314, 79.85975, 80.30109,
    80.10844, 79.97185, 80.49149, 81.30732, 81.44389, 78.77293, 72.48772,
    73.1268, 70.63235, 67.35307, 68.37753, 68.09903, 67.43285, 66.94666,
    66.46853, 66.44505,
  76.94654, 78.49357, 79.03192, 78.72236, 78.00905, 78.05085, 78.29025,
    78.56119, 78.6127, 78.95976, 79.67343, 80.17328, 80.66796, 81.14526,
    80.84134, 80.64712, 80.91788, 77.75621, 73.73655, 72.36694, 71.15222,
    70.46969, 68.47654, 67.67641, 67.99095, 68.03099, 67.35482, 66.80042,
    66.50986, 66.47343,
  78.48167, 77.1544, 77.14391, 77.38065, 77.44586, 77.35592, 77.85371,
    78.28589, 78.22501, 78.28065, 78.86546, 80.04002, 81.47451, 82.05897,
    82.16718, 82.46739, 82.99269, 81.81539, 77.70205, 74.74057, 71.66161,
    71.21432, 69.6511, 68.46719, 68.43736, 68.26861, 67.28073, 66.43498,
    66.34946, 66.4505,
  85.33881, 81.28326, 78.46271, 77.72536, 77.70952, 77.3671, 77.49887,
    77.96459, 78.39877, 77.82732, 77.96505, 78.86295, 80.07261, 81.12595,
    81.94064, 82.99672, 84.38916, 85.60142, 86.07668, 82.34394, 76.07806,
    72.51235, 70.79466, 69.93288, 69.28513, 68.70455, 67.56193, 66.52308,
    66.30689, 66.40471,
  94.70171, 89.67217, 82.70218, 77.48769, 78.70696, 77.92312, 77.98286,
    78.21275, 77.61618, 77.57436, 77.57925, 76.62824, 74.74962, 74.33907,
    75.00304, 78.10782, 83.17754, 85.70946, 87.42044, 88.37104, 83.59703,
    76.36763, 72.32466, 71.69628, 70.28337, 69.38681, 68.26887, 66.82746,
    66.41171, 66.43043,
  93.91859, 90.20726, 84.19389, 79.53713, 80.52539, 80.09021, 80.03825,
    79.82825, 80.01682, 80.54143, 80.41074, 79.39986, 78.92854, 75.91071,
    73.38456, 72.85554, 74.39931, 77.52608, 79.51138, 80.85907, 81.18118,
    78.48739, 74.4417, 72.9595, 71.32395, 69.8746, 68.61401, 67.09489,
    66.37714, 66.51123,
  93.43017, 90.47118, 85.23375, 81.32021, 82.46225, 82.41222, 82.62397,
    82.59844, 82.71667, 82.46288, 81.22559, 80.08973, 80.72158, 79.96362,
    77.79295, 77.00477, 76.80336, 77.2674, 77.68359, 76.57547, 76.38353,
    77.01632, 76.26159, 74.25158, 72.73346, 70.58321, 68.91801, 67.17619,
    66.35189, 66.40883,
  91.79297, 89.85672, 84.73866, 82.36252, 83.65614, 83.95412, 84.51431,
    84.78796, 85.17139, 85.46577, 85.10599, 83.75572, 82.98804, 82.1227,
    80.94666, 80.13802, 79.51888, 79.44993, 79.19303, 77.76196, 75.78304,
    75.04462, 77.08122, 75.41732, 74.48125, 71.90385, 69.7864, 67.87037,
    66.45444, 66.35055,
  90.20103, 88.46745, 83.49482, 81.37029, 82.5625, 83.02527, 83.98359,
    84.95508, 86.45665, 87.69984, 88.1254, 88.04136, 87.73018, 87.424,
    86.98418, 86.42632, 85.21107, 84.10676, 82.72444, 81.21948, 78.95136,
    76.78535, 77.51675, 76.21032, 76.15907, 73.97188, 71.24053, 68.91287,
    67.43242, 66.61314,
  87.84447, 85.75072, 81.71017, 79.88522, 80.63815, 81.1176, 82.32719,
    84.23267, 86.72547, 88.27518, 89.13002, 90.50851, 92.05594, 92.73816,
    92.13245, 92.01727, 91.67454, 90.4744, 88.44505, 86.49171, 84.84657,
    82.23903, 79.33821, 78.05627, 77.77987, 76.6608, 74.1167, 70.467,
    68.79957, 67.47495,
  86.5531, 83.54859, 79.48981, 76.97971, 77.64439, 78.11121, 80.19202,
    82.87611, 85.60556, 86.47463, 87.21649, 88.78244, 91.19057, 92.40664,
    92.06956, 92.09991, 91.81299, 90.88275, 88.86982, 87.83305, 86.13221,
    83.86419, 80.74147, 78.47823, 78.3706, 77.12572, 75.38638, 71.62459,
    69.0427, 67.82936,
  86.9698, 83.71064, 80.20561, 76.51576, 75.99251, 75.66612, 78.17836,
    82.30015, 85.11056, 85.41489, 87.12116, 88.89944, 91.10442, 92.21652,
    92.12859, 92.00309, 90.53443, 89.18053, 88.05164, 87.35587, 85.74763,
    83.84408, 81.34524, 79.58094, 79.36335, 77.97484, 76.32927, 72.81268,
    68.91562, 67.37828,
  88.77711, 86.5313, 81.243, 76.89388, 76.54268, 75.34594, 76.50342,
    78.57496, 79.97952, 80.05159, 82.13484, 84.93423, 88.07787, 89.26487,
    88.1496, 87.82437, 86.66546, 85.8137, 86.15925, 85.32793, 83.85465,
    82.32829, 80.40009, 79.30258, 79.1163, 78.08491, 77.22922, 74.88435,
    70.37752, 67.47369,
  86.14479, 84.47618, 80.49611, 77.46545, 78.27602, 77.72939, 76.90585,
    76.47251, 75.87083, 75.6252, 76.15354, 78.04836, 80.87238, 82.08365,
    81.91453, 81.69839, 80.41561, 79.53947, 79.65959, 80.95752, 80.25259,
    79.00128, 77.0308, 75.96389, 76.03368, 75.10364, 74.30611, 73.91685,
    71.99063, 68.33794,
  73.12401, 74.21187, 75.27094, 75.60041, 76.44923, 78.05373, 76.49178,
    73.20314, 71.97403, 72.17793, 71.80877, 71.47984, 71.91002, 72.60416,
    72.74373, 72.86746, 72.27426, 71.49834, 71.24789, 71.38311, 72.09072,
    72.94697, 72.90552, 72.10677, 72.01595, 71.78362, 71.16245, 69.86906,
    68.95875, 68.14129,
  69.96175, 70.4297, 71.03398, 70.99084, 71.74627, 73.30019, 73.55435,
    71.20507, 69.79602, 70.2377, 70.27956, 70.23912, 70.04438, 69.73643,
    69.4983, 69.4571, 68.93041, 67.96358, 67.75112, 67.70954, 67.51707,
    68.14175, 69.04801, 69.33629, 69.19798, 69.22083, 68.83562, 68.02066,
    67.35506, 66.69054,
  77.73868, 78.14349, 78.1629, 78.16218, 77.80656, 77.5611, 77.37434,
    77.24017, 77.38271, 77.89368, 78.85493, 79.62283, 79.4511, 80.091,
    80.4994, 80.07082, 79.21706, 77.88774, 75.78049, 73.28984, 70.43504,
    67.20073, 65.61513, 65.53632, 64.40924, 60.62141, 58.39507, 60.26241,
    56.25745, 54.07163,
  81.79446, 82.54411, 82.45088, 82.91607, 82.62318, 82.30593, 82.0251,
    81.41678, 80.76602, 80.21105, 79.9852, 80.33102, 80.94656, 81.06821,
    81.50646, 82.61804, 83.6056, 83.34516, 82.28671, 81.16837, 80.11491,
    79.26687, 78.74892, 78.97183, 79.06155, 71.08592, 56.64867, 58.54024,
    56.24286, 54.4516,
  82.15247, 83.08079, 83.87012, 84.64462, 85.21367, 85.78369, 86.13559,
    86.21602, 85.94072, 85.07607, 83.72353, 82.46748, 81.21152, 80.31734,
    79.49959, 78.2457, 78.6673, 80.77524, 82.57504, 81.8332, 81.31596,
    80.90628, 80.64524, 80.56254, 79.93447, 78.10403, 70.48975, 59.61968,
    55.35048, 54.54384,
  82.42847, 83.33026, 84.04874, 84.81615, 85.47282, 86.17006, 86.81194,
    87.16874, 87.29245, 87.1157, 87.11698, 87.7151, 87.75826, 86.89783,
    85.20625, 83.10412, 79.99413, 78.63422, 80.97463, 82.15768, 81.46278,
    80.49104, 80.11694, 80.51876, 79.93466, 78.7564, 77.79619, 75.34712,
    62.35921, 55.66785,
  82.56982, 83.53478, 84.27736, 84.91755, 85.35109, 86.10341, 87.03539,
    87.42881, 87.26904, 86.9211, 87.07922, 88.2348, 88.93723, 88.23494,
    87.4339, 86.7888, 85.29951, 83.53969, 82.73541, 82.24641, 80.96883,
    72.26633, 72.68766, 77.5623, 79.59019, 79.00801, 78.7696, 79.31479,
    78.98208, 65.34341,
  82.50758, 83.73949, 84.61676, 85.2753, 85.63248, 86.54893, 87.86494,
    88.52509, 88.4502, 88.21585, 88.25081, 89.09858, 89.7678, 89.16773,
    89.01501, 88.32365, 86.18472, 84.421, 82.41624, 81.56662, 79.86234,
    68.93134, 72.79543, 74.44469, 77.86063, 79.13312, 79.41834, 80.10696,
    78.96919, 58.6674,
  82.67963, 83.77819, 84.62917, 85.34245, 85.88465, 87.00125, 88.54826,
    89.60357, 89.72236, 89.4156, 89.22592, 88.53596, 82.05115, 82.09563,
    81.83231, 81.55933, 82.43523, 81.87896, 79.06421, 78.52114, 75.18788,
    72.43589, 73.89468, 75.87482, 76.89082, 77.53556, 79.30102, 79.53711,
    75.79562, 52.95117,
  83.69509, 84.42388, 85.18607, 85.87482, 86.32484, 87.37425, 88.48641,
    88.10271, 83.17404, 85.2811, 84.66248, 83.12869, 82.04659, 81.46996,
    81.08186, 80.8193, 80.17191, 78.35034, 75.96751, 74.4407, 73.8465,
    74.45366, 76.24377, 77.87, 78.38551, 78.90015, 79.33408, 78.78777,
    66.30493, 53.18197,
  86.12093, 86.45796, 86.72376, 87.03569, 87.20172, 87.36836, 83.31517,
    81.30315, 82.03947, 81.62728, 82.2182, 82.7507, 83.29183, 85.85716,
    87.2427, 85.27793, 85.18513, 85.23541, 83.92604, 80.45902, 77.28435,
    77.10564, 78.23736, 78.30815, 78.72339, 79.4786, 79.2078, 74.42529,
    53.50599, 54.09338,
  90.12919, 90.13577, 89.72477, 89.51636, 89.22426, 88.07288, 84.00996,
    87.19952, 83.68539, 81.22157, 78.65479, 78.46629, 77.88673, 77.63985,
    78.05688, 79.82335, 81.24625, 81.80215, 82.43378, 83.24844, 82.17699,
    80.47474, 78.05194, 75.9557, 78.5789, 79.24437, 78.25247, 59.80201,
    53.28367, 53.11728,
  94.77587, 94.4326, 95.21788, 93.66449, 93.01881, 90.46323, 88.73803,
    87.65578, 87.35111, 87.256, 80.24809, 73.22144, 72.43871, 71.16072,
    70.1571, 70.23782, 70.35232, 70.701, 72.21042, 75.5293, 80.71957,
    80.70524, 78.27416, 78.28025, 78.71725, 78.2373, 61.82265, 53.66912,
    54.31422, 53.25558,
  98.70989, 97.51594, 100.1635, 100.5812, 98.54986, 95.1561, 91.87956,
    88.56038, 86.78738, 86.87774, 85.69904, 84.33183, 81.98464, 80.06503,
    77.00681, 72.82969, 72.01263, 70.19149, 69.21292, 70.14466, 74.37934,
    76.60002, 75.33609, 78.78896, 78.82462, 73.86359, 54.05036, 58.36686,
    54.94591, 53.82389,
  90.95358, 93.25622, 95.58646, 97.51382, 98.62222, 97.60516, 91.65288,
    87.32348, 88.8679, 87.34489, 86.50755, 85.58795, 85.44598, 85.38739,
    84.62939, 77.99503, 79.65014, 78.63584, 76.00803, 72.81384, 74.19804,
    75.34135, 71.59438, 65.90424, 65.21992, 62.84054, 55.00997, 56.66592,
    56.11576, 54.63136,
  85.20388, 86.46429, 86.9817, 86.67909, 86.77779, 87.55717, 89.07832,
    89.52419, 87.48817, 87.52205, 86.8634, 85.36001, 85.10278, 85.0267,
    83.94704, 83.22595, 82.92908, 82.56763, 82.34786, 81.0997, 77.04007,
    73.19082, 65.02197, 57.84481, 54.14666, 54.65107, 54.21512, 53.79278,
    54.11614, 54.01164,
  85.42357, 86.45811, 86.69025, 86.23705, 85.64126, 85.61135, 86.95443,
    86.88631, 84.38345, 82.82997, 81.71355, 80.72673, 83.071, 82.81077,
    84.58238, 84.58956, 83.00959, 81.66703, 78.8573, 74.87672, 67.74102,
    63.69962, 57.88054, 55.38132, 55.95352, 55.4589, 54.64333, 53.98773,
    53.50192, 53.3555,
  80.52947, 84.02724, 85.8024, 86.43727, 87.01469, 88.23513, 89.20731,
    89.43415, 88.51772, 84.77237, 83.08208, 81.43725, 80.8158, 82.28795,
    79.53709, 77.91519, 78.54055, 73.41718, 68.90741, 64.97321, 61.52264,
    59.83992, 56.39526, 55.25964, 55.65194, 55.51073, 54.46836, 53.91408,
    53.59964, 53.40482,
  77.40044, 77.50896, 78.62972, 80.22298, 81.8426, 83.4303, 85.69354,
    88.81927, 89.52377, 88.4734, 86.26651, 87.77246, 88.79517, 88.36964,
    83.9413, 81.94987, 78.86462, 76.01701, 71.89213, 67.68822, 62.54276,
    60.78476, 57.5018, 55.72244, 55.68805, 55.4891, 54.30437, 53.48233,
    53.38651, 53.36464,
  82.38704, 79.82697, 77.73156, 77.61118, 78.18427, 79.22219, 80.88769,
    82.99686, 84.77366, 85.18837, 87.11657, 88.49486, 89.17546, 88.84982,
    88.04564, 88.54725, 88.64423, 86.66911, 81.73457, 74.78737, 66.38293,
    61.82843, 58.88612, 57.33857, 56.00033, 55.32132, 54.43784, 53.41815,
    53.25888, 53.25589,
  96.18222, 90.2222, 81.37074, 76.25243, 77.41355, 77.04379, 77.91108,
    78.83301, 78.78799, 79.40496, 80.46114, 79.59396, 77.34589, 77.08308,
    77.22456, 79.88003, 85.4034, 89.55638, 88.4439, 83.37698, 74.34452,
    65.57016, 60.58418, 58.92596, 57.10066, 55.96965, 54.95399, 53.68119,
    53.29605, 53.31371,
  97.10005, 92.96696, 84.06245, 78.84268, 79.55221, 79.22603, 79.54678,
    79.85128, 80.37335, 81.21352, 81.16687, 79.29763, 78.45639, 75.00337,
    71.91847, 71.00414, 72.82027, 76.40318, 77.31652, 76.40427, 73.429,
    68.31516, 63.06478, 60.41094, 58.49327, 56.55436, 55.28272, 53.83897,
    53.26701, 53.32372,
  98.22523, 95.94233, 87.54314, 82.88236, 83.29107, 82.70026, 82.74846,
    82.73047, 82.96072, 82.92488, 81.33035, 79.97956, 80.76517, 79.33037,
    76.93137, 75.49738, 74.75845, 74.6212, 74.04608, 71.06314, 68.90751,
    67.54462, 65.07113, 62.53926, 60.02407, 57.3574, 55.41463, 53.97646,
    53.23502, 53.29724,
  98.85527, 97.64033, 90.99104, 87.63198, 88.75662, 87.9834, 87.98179,
    87.83258, 88.27343, 87.77001, 85.43926, 83.3875, 82.76518, 81.53188,
    79.82645, 78.40423, 76.5871, 75.45799, 74.41341, 72.44815, 70.0559,
    66.94947, 65.25391, 64.12747, 62.03206, 58.53055, 56.2718, 54.64825,
    53.44665, 53.23074,
  99.74713, 98.99942, 92.21433, 89.47807, 91.81964, 92.29414, 92.47303,
    92.57447, 93.98428, 93.7448, 91.91674, 91.83037, 91.01012, 89.30903,
    87.02361, 84.78233, 81.79024, 78.49557, 75.93623, 73.38192, 70.77855,
    67.49368, 64.83949, 64.13705, 63.99441, 61.0359, 57.71611, 55.82407,
    54.40752, 53.42627,
  100.1446, 98.4445, 92.10001, 89.72412, 90.88725, 90.70314, 92.13896,
    94.23621, 98.31435, 98.69344, 97.31357, 99.13203, 100.7707, 100.1483,
    97.48444, 94.72547, 90.85688, 86.28484, 82.19657, 78.31033, 74.1853,
    70.4024, 67.0415, 65.6096, 65.53519, 64.56243, 61.38805, 57.48668,
    55.75173, 54.24937,
  101.2383, 96.0169, 88.82422, 85.43918, 85.45367, 85.08829, 87.93864,
    93.22051, 98.48328, 97.28578, 95.32189, 96.95786, 99.13498, 99.54625,
    97.59755, 95.37402, 91.71838, 88.04529, 85.32012, 82.24081, 77.66887,
    73.14233, 68.7216, 66.12687, 66.12029, 65.39436, 63.60924, 59.33349,
    56.36441, 54.8682,
  100.0906, 95.42296, 89.11443, 84.70554, 83.21445, 81.98828, 85.09745,
    90.67104, 94.23854, 92.674, 93.13026, 94.23727, 96.2662, 96.83991,
    94.81512, 92.17619, 89.19468, 86.16157, 84.18427, 82.18092, 78.67615,
    74.74996, 70.61369, 68.08061, 67.53341, 66.13687, 64.68413, 60.61371,
    56.01853, 54.36108,
  95.45728, 91.8497, 86.06063, 82.07613, 81.00209, 78.69342, 80.0223,
    82.38461, 84.01266, 83.4085, 84.87469, 86.91761, 89.164, 89.74648,
    88.65526, 86.71382, 83.81701, 81.59143, 80.69305, 79.07656, 75.85889,
    73.57507, 71.03609, 69.1686, 68.8192, 67.92992, 67.04107, 63.86912,
    57.67271, 54.06353,
  85.60069, 83.95147, 80.82354, 77.71382, 78.42047, 77.02979, 75.44275,
    74.3093, 72.74596, 72.4338, 72.86648, 74.4105, 76.82674, 77.81721,
    77.02148, 76.45246, 74.21516, 72.66118, 72.76307, 72.59747, 70.73228,
    68.32507, 65.66107, 64.55893, 64.74393, 64.25885, 63.50381, 62.89563,
    60.55614, 55.41391,
  68.04709, 69.121, 69.61021, 69.61604, 70.71254, 72.38715, 69.75646,
    65.21334, 63.5834, 63.887, 63.33806, 62.98602, 62.97935, 63.30324,
    63.32775, 63.1627, 62.62487, 61.63043, 61.02629, 60.98936, 60.8756,
    61.15992, 60.84519, 59.83804, 60.04758, 59.99073, 59.01506, 57.51211,
    56.70039, 55.34241,
  60.37135, 61.04205, 61.36289, 60.73205, 61.34357, 63.278, 63.81852,
    60.17804, 58.2783, 59.13653, 59.65165, 59.57803, 59.42057, 58.85796,
    58.14429, 57.95736, 57.07661, 55.69871, 55.54966, 55.43385, 55.00727,
    55.5694, 56.41828, 56.87059, 56.78215, 56.95767, 56.58881, 55.34683,
    54.37214, 53.45412,
  66.87151, 66.67416, 66.40607, 66.481, 66.37776, 66.42002, 66.67276,
    66.97605, 67.35535, 67.98764, 69.18893, 68.74493, 65.589, 64.89072,
    63.96694, 62.07902, 60.52862, 59.44057, 58.35406, 57.76809, 56.56477,
    54.39806, 54.28773, 55.9236, 56.52562, 54.15192, 54.9685, 56.52084,
    46.70355, 42.84808,
  73.40699, 73.0753, 71.63972, 71.70576, 70.80174, 70.26679, 70.36472,
    70.61153, 71.06484, 71.72113, 72.89151, 74.37203, 75.12917, 73.84141,
    72.40461, 72.07853, 70.76839, 70.57888, 70.52433, 70.36207, 69.30959,
    68.22882, 67.61764, 69.5966, 70.77922, 60.89978, 50.62096, 53.50564,
    46.75787, 43.7003,
  76.22503, 76.5282, 76.09048, 75.48266, 74.84566, 74.12316, 73.17677,
    72.54128, 72.0733, 71.65257, 71.57577, 72.10632, 72.96498, 74.29662,
    74.92746, 73.20135, 73.20528, 74.53312, 76.10902, 78.47935, 82.64649,
    83.123, 83.22972, 83.35461, 79.97607, 70.93674, 61.31862, 53.0232,
    45.78497, 43.9991,
  79.94849, 80.55021, 81.08921, 81.56392, 81.27155, 81.09406, 80.83156,
    79.95998, 79.20898, 78.31461, 77.51534, 77.50288, 76.45056, 75.03329,
    76.48763, 76.40874, 73.16617, 71.38357, 74.74409, 79.1273, 82.95603,
    82.88657, 78.86657, 82.57246, 79.62687, 76.32793, 72.24969, 62.32914,
    50.57963, 44.20515,
  82.55186, 82.33742, 82.11833, 81.69422, 81.20358, 81.0308, 81.10232,
    80.80761, 80.50041, 80.18417, 80.26466, 81.11892, 81.78233, 81.89235,
    82.1208, 82.50319, 81.90583, 76.51975, 76.33978, 80.15338, 76.98996,
    67.24627, 68.48637, 74.42717, 79.25074, 79.72824, 78.49449, 81.16148,
    77.07702, 53.33879,
  82.73335, 82.91113, 82.72183, 82.29681, 81.48986, 81.44497, 82.13792,
    81.84634, 81.11096, 80.63415, 80.82402, 81.82236, 82.81022, 82.96582,
    83.83165, 84.59399, 83.8021, 82.31363, 81.21494, 79.27783, 70.77531,
    61.82085, 66.60905, 70.28415, 75.18172, 77.40202, 79.50053, 82.36844,
    80.85388, 48.04313,
  81.32975, 83.03619, 83.07066, 82.7408, 82.09992, 82.35334, 83.2165,
    83.16658, 82.53187, 81.97539, 81.78822, 81.38409, 75.47948, 77.10372,
    78.92617, 80.33829, 80.16006, 76.44008, 71.23435, 71.18736, 67.65819,
    65.3865, 68.04075, 71.89155, 73.10478, 70.94707, 74.27273, 78.94899,
    65.87002, 41.50449,
  82.11504, 83.10542, 83.26559, 83.22125, 82.93813, 83.28144, 83.95341,
    83.09264, 82.22945, 82.1778, 81.39592, 79.04794, 77.34146, 77.13934,
    76.91891, 77.54573, 78.58763, 76.56014, 71.94362, 70.144, 69.33916,
    70.82138, 74.35266, 76.00371, 73.90821, 74.92023, 79.85297, 75.17842,
    57.64012, 42.64125,
  84.1712, 84.03853, 83.72487, 83.23852, 82.42863, 82.36716, 82.10292,
    82.82529, 83.39366, 83.5173, 83.67525, 83.72601, 83.99429, 85.3048,
    86.0472, 84.96499, 85.23878, 85.58761, 84.44742, 78.2468, 73.92992,
    76.21487, 80.59303, 79.59376, 76.14594, 81.90193, 80.20301, 65.65909,
    43.82449, 42.81479,
  85.65817, 86.21333, 85.21658, 84.98162, 83.96577, 82.18914, 78.55714,
    81.62628, 82.04343, 82.76584, 83.16399, 83.42796, 83.08388, 82.2971,
    81.01525, 84.3649, 85.02401, 84.8174, 83.05891, 83.77656, 84.28305,
    79.24715, 73.70714, 68.40595, 73.80396, 80.92384, 70.22582, 50.98973,
    42.08676, 41.05276,
  86.19695, 86.00673, 87.30319, 85.53241, 85.87551, 83.6949, 82.47742,
    81.98355, 82.64834, 83.61091, 80.34489, 66.53635, 63.12896, 63.05081,
    62.59724, 63.90758, 65.30582, 65.96775, 67.24717, 72.08609, 80.55999,
    77.0357, 68.19724, 67.99587, 72.34933, 67.48676, 51.20313, 43.00707,
    43.02807, 41.30089,
  91.66879, 89.73187, 91.56821, 92.05653, 89.2922, 86.70281, 84.3194, 81.661,
    80.10192, 80.09026, 78.30306, 76.78263, 77.01552, 74.87, 65.57851,
    64.94495, 63.29884, 62.40322, 62.25864, 64.90809, 72.1441, 73.55352,
    66.65305, 73.77802, 76.43074, 62.55081, 43.78125, 47.59572, 44.23737,
    42.30767,
  89.36157, 90.99651, 92.57267, 93.38536, 92.82886, 90.58459, 84.344,
    80.86396, 82.41283, 81.53379, 81.87772, 81.6787, 82.79957, 83.17381,
    81.38184, 70.94135, 70.12462, 69.00221, 66.92039, 67.63242, 70.06384,
    68.5817, 63.24505, 58.4917, 57.32479, 53.1743, 44.76824, 46.37936,
    45.80621, 43.44236,
  82.16991, 82.69135, 83.18056, 82.12029, 81.85361, 82.3849, 83.58635,
    83.80562, 81.90871, 82.69571, 83.35368, 83.10648, 84.44746, 84.79043,
    83.07362, 81.29755, 78.15573, 81.73333, 82.56219, 75.86462, 69.23867,
    64.21763, 55.95295, 48.78003, 45.23244, 44.92842, 43.49579, 42.70517,
    43.07726, 42.62881,
  85.13036, 85.25323, 83.90601, 82.59448, 81.84781, 82.4681, 84.28976,
    84.33806, 82.34074, 82.21128, 82.04794, 81.47965, 81.8942, 82.81743,
    82.50211, 81.14112, 80.58749, 78.11475, 77.62994, 71.53359, 59.20227,
    55.25334, 48.75373, 46.40486, 46.4656, 45.45596, 44.01354, 42.96406,
    42.06784, 41.65261,
  85.36301, 85.956, 85.78054, 84.90173, 84.21644, 84.68321, 85.26015,
    84.58833, 83.19704, 79.89639, 77.90107, 74.71382, 72.69093, 75.74229,
    73.3988, 72.15005, 73.04414, 69.18335, 66.74613, 60.71513, 52.7943,
    52.08204, 47.29229, 45.80738, 45.99671, 45.33153, 43.54766, 42.86636,
    42.31662, 41.7052,
  79.36035, 79.31664, 80.96238, 83.59568, 83.90257, 83.63494, 84.09375,
    85.11785, 84.79203, 83.75391, 82.5137, 83.09759, 84.38983, 83.53401,
    77.18153, 74.18536, 70.70628, 68.93359, 67.31583, 62.23634, 52.88329,
    52.65955, 48.66391, 46.10921, 45.6405, 45.27229, 43.23257, 41.78487,
    41.73654, 41.5812,
  77.83842, 77.12595, 75.3868, 76.67667, 78.1761, 80.30375, 82.78902,
    84.12377, 84.73884, 84.3391, 84.8922, 85.62559, 85.68592, 85.77964,
    84.97685, 84.88645, 83.02664, 81.36919, 77.22771, 68.27331, 55.50386,
    52.08654, 49.0878, 47.6363, 45.29288, 44.18723, 43.33976, 41.58363,
    41.37115, 41.28047,
  90.01038, 83.43935, 74.78564, 70.70923, 72.24795, 72.37885, 73.93484,
    75.86595, 76.40788, 78.45263, 81.72515, 79.83691, 74.68192, 76.42545,
    77.13731, 80.63694, 87.80574, 90.22943, 89.80016, 81.80288, 66.45588,
    56.17618, 50.86605, 48.38953, 45.78616, 44.15381, 43.23164, 41.88062,
    41.36821, 41.29421,
  89.05056, 83.71255, 75.80535, 70.75673, 71.41801, 71.48663, 72.09032,
    73.01561, 74.85374, 77.82545, 77.18294, 70.96798, 70.50311, 68.3677,
    65.89218, 64.96347, 68.47925, 74.60339, 77.31899, 76.08802, 70.37113,
    62.26442, 54.74669, 50.61512, 47.79425, 44.84467, 43.39399, 42.06424,
    41.37182, 41.34956,
  90.81027, 86.25833, 77.96091, 73.30975, 72.82809, 72.18787, 72.3329,
    72.94595, 74.42994, 75.50758, 71.82419, 67.8912, 70.60551, 69.65045,
    67.06874, 65.08843, 65.00294, 65.85738, 66.84077, 65.41112, 64.41288,
    64.12244, 60.34435, 55.0104, 50.18272, 46.04044, 43.53442, 42.17164,
    41.41018, 41.34783,
  95.63418, 91.99638, 84.47204, 80.87986, 80.55159, 78.37575, 77.85862,
    77.38273, 78.93202, 78.02554, 72.01751, 69.17679, 70.18552, 69.28896,
    67.52869, 66.46709, 64.54079, 63.50204, 63.44754, 63.00408, 62.51464,
    61.21445, 60.87465, 59.88628, 54.94012, 47.92471, 44.51436, 43.15936,
    41.69562, 41.30444,
  98.15468, 97.09773, 90.14211, 87.32166, 89.20126, 88.63721, 86.66219,
    84.64137, 85.27663, 82.90832, 77.39081, 77.63326, 77.29062, 76.10896,
    73.72348, 72.23024, 69.50822, 65.26333, 62.60232, 61.1666, 60.16786,
    58.44627, 57.11125, 58.27599, 58.80372, 52.81807, 47.05919, 45.18724,
    43.20848, 41.53441,
  97.89889, 96.56682, 92.50568, 90.40871, 90.39793, 88.85226, 88.97953,
    89.81443, 93.54745, 90.68597, 85.36016, 87.8603, 89.29491, 88.93311,
    86.00298, 83.30225, 79.66243, 74.63374, 68.9644, 64.99791, 62.34377,
    59.89785, 57.66096, 57.07873, 58.15216, 58.30117, 53.56112, 47.69767,
    45.40082, 42.75687,
  97.43149, 94.52816, 86.79419, 83.1498, 82.3427, 81.0649, 83.60914,
    89.70187, 94.6825, 91.0267, 85.09967, 87.38537, 89.10069, 89.69421,
    87.89613, 86.3924, 83.29359, 79.91367, 75.94621, 71.45692, 67.32486,
    63.55236, 59.8618, 57.23972, 57.61608, 58.28926, 57.34999, 51.32596,
    47.12955, 44.32487,
  95.59586, 93.21906, 89.04921, 83.38922, 80.07487, 78.30733, 82.69864,
    89.61758, 92.08198, 86.82118, 86.18169, 87.25021, 88.79506, 88.27739,
    85.78849, 84.58817, 83.16933, 80.92754, 78.83747, 76.16111, 73.44318,
    70.14518, 65.89264, 62.46264, 61.72895, 60.42638, 59.63817, 53.97572,
    45.76462, 43.27691,
  92.51836, 90.39478, 86.16436, 81.67935, 79.30676, 76.2662, 79.02421,
    82.00976, 82.03872, 79.93862, 81.81615, 83.59736, 84.55768, 83.77374,
    82.40008, 80.65884, 78.81672, 77.70865, 76.79401, 75.11268, 73.30615,
    72.89922, 71.82558, 69.25301, 68.34492, 67.37971, 67.61637, 62.84985,
    49.53216, 42.1904,
  85.64747, 84.9871, 82.96933, 82.0234, 82.89426, 81.22104, 78.96152,
    75.68832, 71.52464, 71.65852, 72.21182, 73.76511, 75.32458, 75.55614,
    74.89912, 73.49547, 71.04887, 70.09451, 70.2441, 70.27074, 67.30138,
    63.13665, 59.93751, 59.4678, 60.86105, 61.58196, 62.16475, 63.27777,
    57.94447, 45.55256,
  70.37307, 71.13691, 71.53902, 72.31801, 75.94069, 79.78485, 75.02136,
    65.79371, 62.71965, 63.42844, 62.4914, 62.04144, 62.24042, 62.42631,
    62.29268, 61.51208, 59.63828, 58.06484, 56.7441, 54.83643, 53.80562,
    53.14416, 51.34705, 50.02304, 51.13102, 52.08072, 51.60081, 49.58043,
    49.02152, 46.19361,
  58.89107, 59.45137, 59.07988, 58.14604, 59.88562, 64.85305, 66.24267,
    57.76197, 53.63906, 56.02359, 57.55737, 58.61395, 58.77614, 57.4706,
    55.42326, 53.82112, 50.53313, 47.332, 46.95692, 46.36643, 44.90901,
    45.48674, 45.97583, 46.12557, 46.48462, 47.45633, 47.41357, 45.23081,
    43.05484, 41.30582,
  51.79374, 51.71765, 51.72526, 51.86572, 51.71323, 51.81242, 52.19237,
    52.69604, 53.4123, 54.5904, 57.1363, 57.14211, 53.13315, 53.7827,
    54.29657, 53.73364, 53.97147, 55.01759, 56.21169, 58.13486, 58.75721,
    57.21792, 58.07742, 61.0733, 63.14267, 62.5443, 67.83218, 69.60841,
    53.81189, 49.49067,
  55.17516, 55.35119, 54.4959, 55.22848, 54.36712, 53.94326, 54.48619,
    55.08757, 55.90007, 56.88635, 58.63681, 61.02748, 62.38475, 60.24068,
    58.82528, 59.68481, 58.66225, 59.90212, 61.85575, 63.35532, 62.98898,
    62.18158, 62.58473, 66.6305, 70.10987, 65.12965, 62.33552, 67.07325,
    54.98304, 50.9502,
  54.17039, 54.51822, 55.26799, 55.89277, 56.25319, 56.53949, 56.57384,
    56.99554, 57.64064, 58.45879, 59.56584, 61.26055, 63.08518, 65.4555,
    66.49554, 64.08781, 64.27689, 65.89917, 67.21304, 69.33863, 72.85979,
    76.50165, 77.91458, 78.28772, 77.71303, 72.69727, 69.47829, 65.23351,
    54.21463, 51.85254,
  56.91003, 57.13821, 58.47077, 59.9238, 61.65506, 63.45611, 63.25208,
    62.49585, 63.22486, 64.1555, 64.71405, 65.76836, 65.63498, 64.88191,
    68.34214, 70.41203, 67.09177, 64.2533, 67.27403, 71.1172, 76.04291,
    76.37383, 74.88431, 80.12979, 80.67635, 78.41309, 73.76739, 65.29388,
    56.02287, 50.53937,
  59.9165, 59.40015, 61.36029, 62.72267, 63.65387, 64.25224, 64.56953,
    64.49973, 66.11594, 67.42933, 68.08048, 70.95889, 72.51238, 73.259,
    74.43587, 76.31575, 73.91597, 67.94964, 69.15701, 74.43363, 74.04387,
    67.07467, 69.04963, 76.1211, 82.62332, 80.12234, 72.24197, 76.39335,
    73.95866, 56.82237,
  61.4665, 63.54361, 67.15646, 70.47208, 70.257, 70.94029, 73.93295,
    74.43521, 73.43208, 74.1888, 76.52602, 82.42739, 86.76868, 87.02228,
    88.04105, 89.33787, 89.22276, 84.14028, 74.60822, 75.26839, 70.42185,
    64.44579, 68.48705, 74.57137, 81.52679, 79.82539, 74.10551, 83.37609,
    78.94377, 54.85214,
  62.12373, 64.45766, 67.59842, 70.41349, 71.21228, 72.93677, 77.02132,
    80.06319, 78.65202, 77.02732, 76.74474, 73.2514, 69.06276, 72.26661,
    75.75537, 78.62274, 81.46966, 77.54762, 69.45248, 71.14042, 69.00276,
    68.05901, 71.69294, 78.21793, 79.20965, 72.33904, 72.54286, 77.51293,
    70.28837, 50.13817,
  62.63608, 64.74117, 68.388, 71.33817, 71.47014, 75.93202, 79.76436,
    71.86344, 66.35249, 67.96638, 68.46736, 68.58796, 69.16048, 73.05135,
    76.30138, 79.33425, 83.45082, 82.56476, 75.9582, 74.11025, 72.91869,
    75.34256, 80.87825, 83.5484, 78.62717, 75.8047, 80.27524, 78.31854,
    66.08824, 50.4497,
  74.36766, 75.22065, 76.84582, 77.16996, 76.41257, 78.62828, 74.71586,
    75.26129, 79.40804, 82.61221, 84.12499, 85.42868, 89.04948, 92.98503,
    94.62499, 92.6403, 93.55538, 94.59136, 94.22273, 91.42641, 84.93321,
    90.42389, 93.60239, 92.37663, 84.32305, 89.62176, 86.81094, 73.14204,
    53.75731, 49.56077,
  88.24155, 89.67388, 89.27602, 89.75865, 88.43797, 86.74693, 76.76386,
    81.44644, 82.44246, 88.70706, 91.40805, 92.73502, 92.46698, 91.16788,
    86.92807, 91.82621, 92.95331, 93.34311, 93.35081, 94.7361, 95.62096,
    93.5004, 91.41611, 81.18812, 80.64685, 83.65696, 75.5684, 58.22886,
    49.31203, 46.8781,
  86.57224, 86.25894, 87.91679, 87.65214, 88.9313, 88.71556, 86.91861,
    88.43484, 89.63882, 90.45386, 81.50179, 64.11581, 63.04107, 63.56168,
    64.6069, 66.51571, 69.78893, 70.79343, 71.98569, 77.859, 91.24366,
    87.5144, 71.14386, 66.62057, 69.95824, 66.84383, 55.78431, 49.74604,
    48.97855, 47.07113,
  91.3825, 89.25581, 92.41412, 92.88654, 90.90204, 89.31077, 84.26299,
    79.19176, 73.50494, 67.93262, 64.53476, 62.36785, 65.1808, 67.08944,
    66.51603, 65.94553, 65.11823, 65.83401, 67.75054, 73.9456, 85.64611,
    83.69968, 67.64811, 73.7884, 75.38346, 63.21667, 50.46792, 52.3615,
    50.46629, 48.21143,
  93.541, 95.28751, 97.09451, 96.99057, 95.93236, 93.25289, 87.27998,
    84.73714, 86.42229, 77.68899, 75.36304, 73.01328, 76.77132, 79.81808,
    77.34177, 69.64307, 71.00875, 71.7756, 76.56116, 85.13387, 82.24464,
    76.46931, 66.81044, 64.6889, 64.05829, 58.35107, 51.41501, 52.24293,
    52.19457, 49.32068,
  85.35384, 86.34602, 87.30336, 86.48489, 86.32529, 87.42279, 89.11113,
    89.33353, 87.034, 87.55672, 88.45605, 87.16296, 88.47485, 89.40659,
    87.94208, 78.53379, 75.36208, 77.97655, 81.37306, 79.97692, 72.21882,
    65.28799, 61.5614, 57.67823, 54.06971, 53.04007, 50.33036, 49.12543,
    49.48662, 48.64516,
  76.67586, 77.30474, 81.56227, 84.13256, 84.4688, 86.32097, 89.42117,
    90.23138, 88.09662, 87.69543, 82.90378, 79.2951, 83.5087, 85.74322,
    84.49862, 84.91205, 80.99599, 80.21003, 82.98204, 78.15947, 59.99827,
    60.77682, 56.95312, 55.45102, 54.86525, 52.73642, 50.72099, 49.35044,
    48.19629, 47.61813,
  75.979, 78.83249, 81.76318, 81.73271, 80.05182, 85.08409, 89.65194,
    89.74181, 83.18658, 79.49628, 80.53372, 75.72096, 72.68495, 78.30444,
    76.13744, 76.18192, 78.6983, 76.90134, 77.98292, 72.14037, 58.46886,
    58.92605, 54.73511, 53.78694, 54.22816, 53.11543, 50.4527, 49.58411,
    48.55594, 47.61872,
  69.56031, 67.60909, 69.81155, 71.92154, 73.73193, 76.0779, 79.94129,
    85.22256, 85.81274, 84.1862, 78.36406, 83.70705, 91.49966, 87.12979,
    77.56792, 75.93149, 73.46523, 72.45549, 76.43868, 73.73358, 57.66387,
    59.66063, 56.35849, 54.01141, 52.88663, 52.64849, 50.09736, 47.80365,
    47.82083, 47.50954,
  63.89331, 64.29768, 63.74643, 66.09674, 68.7421, 73.38771, 76.08376,
    76.86188, 80.29822, 79.61837, 88.92566, 92.27589, 92.66521, 91.31725,
    89.53574, 84.39684, 76.61758, 77.36786, 83.26744, 73.80917, 59.19855,
    57.67656, 55.95409, 54.8298, 51.93263, 50.66071, 49.87747, 47.54056,
    47.33841, 47.11706,
  70.30296, 66.29937, 61.29234, 59.49705, 61.37098, 62.45554, 64.69579,
    67.23838, 67.76452, 71.96034, 80.02783, 79.96301, 71.4443, 73.62851,
    75.70218, 79.39495, 86.78452, 94.43436, 96.51239, 88.97688, 69.96368,
    60.21444, 56.35437, 54.34533, 51.30935, 49.73372, 49.1229, 47.7947,
    47.27517, 47.07944,
  68.58678, 65.67485, 60.56808, 58.08652, 59.24768, 60.26772, 61.50112,
    63.2457, 66.90628, 74.90454, 77.5375, 69.13348, 68.62247, 67.48971,
    66.39307, 66.71786, 71.14524, 78.01357, 82.30891, 83.2811, 76.6646,
    67.58231, 59.34287, 56.03441, 53.52187, 50.48724, 49.19539, 47.82903,
    47.27711, 47.10316,
  65.17269, 63.17607, 58.42964, 56.66678, 56.81441, 57.61189, 58.76071,
    60.58905, 64.75957, 70.30131, 67.49949, 62.27225, 67.07549, 67.13593,
    65.6283, 64.4286, 66.07433, 67.74649, 68.65057, 68.52669, 69.5914,
    71.46474, 67.13962, 61.56005, 56.33344, 51.85507, 49.06213, 47.82719,
    47.3158, 47.13031,
  65.70734, 61.5017, 58.69456, 57.87817, 58.48075, 57.43764, 58.55711,
    59.73283, 65.16546, 67.54533, 60.12611, 56.36602, 59.78906, 61.00984,
    61.29394, 62.3194, 62.51388, 63.30231, 65.175, 65.83297, 66.11939,
    67.3097, 69.51399, 68.82413, 61.40466, 53.09237, 49.17655, 48.62907,
    47.60823, 47.16718,
  68.52605, 67.86117, 63.50786, 61.6785, 65.8513, 67.60712, 66.62652,
    64.61672, 66.69329, 64.80448, 57.43305, 58.41465, 60.49211, 62.25902,
    62.27556, 64.17927, 64.826, 62.19262, 61.46383, 61.39145, 60.66387,
    60.67942, 60.97862, 63.82138, 65.769, 58.40858, 51.6501, 50.65796,
    49.13986, 47.39822,
  72.69479, 72.00935, 70.28217, 69.10456, 70.95614, 70.64388, 72.93713,
    74.3647, 77.97848, 71.2656, 62.27773, 64.83208, 66.90571, 69.31016,
    69.46276, 70.03396, 70.73159, 68.87052, 65.12381, 63.23564, 61.42203,
    60.34056, 60.04833, 60.18669, 62.66719, 65.36886, 60.17817, 52.83807,
    51.31203, 48.45914,
  77.9971, 74.36076, 67.15289, 65.45536, 67.97522, 68.66334, 69.41014,
    73.41665, 80.08241, 75.56726, 65.84685, 67.51588, 68.51322, 70.04804,
    71.01686, 72.9808, 73.61248, 73.61019, 70.92328, 67.47394, 65.14237,
    63.73924, 62.23562, 60.75868, 61.12606, 64.58533, 65.89656, 59.06051,
    54.97974, 51.06946,
  82.38863, 80.96205, 75.99222, 69.97799, 68.57032, 68.41554, 73.5321,
    79.16615, 78.4786, 73.16477, 71.87038, 71.3744, 71.58444, 71.39664,
    70.7366, 73.1132, 75.65404, 76.81403, 76.28403, 73.69775, 71.67996,
    70.18338, 66.76759, 63.68136, 63.58133, 64.49731, 66.86829, 61.81804,
    53.19195, 50.07337,
  83.01024, 79.44835, 73.94299, 69.64814, 68.88223, 66.7041, 71.72673,
    74.27539, 70.82487, 69.24075, 72.05589, 72.32963, 71.74037, 71.41653,
    72.32828, 73.9233, 76.244, 78.90001, 80.18642, 79.33676, 78.61198,
    81.10171, 81.83311, 78.14125, 75.76028, 74.90759, 77.25504, 72.54902,
    56.81107, 47.86354,
  79.36269, 74.80367, 75.08583, 75.04843, 77.95187, 76.57289, 75.06183,
    70.79163, 64.40717, 66.50255, 68.00579, 68.72227, 69.15173, 69.84619,
    71.84112, 72.78342, 72.63931, 74.31518, 76.84032, 78.54109, 75.79781,
    71.66279, 69.42385, 69.49877, 70.38165, 71.49093, 73.07695, 76.05988,
    69.58621, 52.5224,
  66.22921, 65.82964, 69.32263, 73.63119, 78.7365, 83.59869, 79.72419,
    67.64468, 63.72451, 65.4097, 65.4202, 66.91584, 68.32509, 69.01247,
    70.34714, 70.50004, 68.89585, 67.30159, 64.17225, 60.52476, 59.31622,
    58.06138, 55.67656, 54.35114, 56.12329, 58.28464, 59.02731, 57.66457,
    57.94854, 53.64118,
  66.35425, 69.65362, 70.27756, 65.68983, 71.15593, 79.60206, 81.72128,
    70.11452, 64.12012, 68.10954, 71.14986, 75.27, 76.21769, 72.25468,
    69.13608, 66.62749, 61.48216, 56.38088, 55.47862, 53.99778, 51.72953,
    51.85548, 51.84401, 51.67709, 52.27514, 53.90892, 54.56005, 52.29745,
    49.37414, 47.10974,
  47.325, 47.92553, 48.44706, 48.99374, 49.44051, 49.98345, 50.58956,
    51.25611, 52.06054, 52.97827, 54.76256, 55.00229, 53.04068, 53.63728,
    53.82369, 53.07783, 52.90369, 53.22635, 53.70554, 54.94711, 55.52166,
    54.81899, 55.51447, 56.74059, 56.94129, 55.77945, 58.65713, 58.434,
    48.36578, 45.22758,
  54.29017, 55.31254, 55.51061, 56.73149, 57.07888, 57.59616, 58.52308,
    59.41477, 60.38572, 61.34227, 62.41346, 63.72672, 64.44312, 62.99651,
    61.90887, 61.709, 60.23582, 60.12712, 60.63879, 61.07957, 60.60504,
    59.73418, 59.82378, 62.40833, 65.81281, 63.21575, 59.20402, 59.97229,
    49.55204, 46.41164,
  57.78033, 59.00466, 60.06907, 61.3396, 62.48637, 63.63519, 64.79543,
    66.14282, 67.44837, 68.54099, 69.46294, 70.5675, 71.58722, 72.91851,
    73.2273, 71.30365, 70.70273, 70.69647, 70.37146, 70.68029, 71.96091,
    73.03905, 72.71829, 72.75231, 73.6385, 70.8679, 65.47697, 59.49048,
    49.97639, 47.45013,
  63.60639, 65.44894, 67.31291, 69.25728, 71.11096, 73.18009, 74.40881,
    75.16067, 76.50931, 77.65685, 77.94146, 78.49052, 78.47615, 77.94542,
    79.67495, 80.17315, 77.04389, 74.01768, 74.14962, 74.7802, 76.96278,
    75.73338, 72.38346, 76.95649, 78.43565, 72.79861, 68.45158, 58.43096,
    50.06189, 46.09722,
  68.90838, 70.08881, 71.96571, 73.80042, 75.1944, 76.42249, 77.5793,
    78.59783, 80.5035, 81.74892, 81.47851, 81.67484, 81.70441, 82.21682,
    82.26001, 81.65573, 78.75854, 74.06053, 73.35903, 77.62823, 77.76646,
    71.13336, 70.96252, 73.62338, 76.61356, 74.20392, 67.5344, 67.57394,
    62.86135, 49.59544,
  76.41068, 79.45574, 82.27275, 85.12778, 85.7016, 86.14202, 88.07616,
    89.28706, 89.12636, 88.6129, 88.2654, 88.49116, 88.30573, 86.94844,
    85.82034, 85.41056, 84.18002, 80.58438, 77.77628, 77.32016, 73.12314,
    68.43625, 69.35847, 70.93465, 73.79987, 71.88781, 69.13981, 75.7053,
    71.58385, 48.24144,
  86.04343, 89.07914, 89.33109, 89.39655, 88.81149, 88.97784, 89.78562,
    89.75668, 88.97649, 88.32539, 87.77137, 86.12433, 81.1255, 80.25163,
    82.6935, 84.57816, 82.70255, 78.39716, 72.19138, 71.48434, 68.93663,
    67.20727, 68.00952, 70.82112, 71.24033, 67.46004, 69.43427, 75.81696,
    65.42693, 45.51194,
  87.20014, 89.47092, 89.72392, 89.84982, 89.35068, 89.27654, 89.78027,
    84.42747, 79.65559, 79.15855, 77.89498, 76.54683, 75.63064, 76.36338,
    77.83084, 78.7506, 78.35635, 75.97527, 71.02708, 69.80899, 68.42301,
    68.34939, 70.50159, 71.76066, 68.40322, 66.394, 71.96467, 70.1917,
    55.68713, 45.82767,
  91.06236, 91.82678, 92.14376, 92.15792, 91.64533, 91.76006, 91.89826,
    91.99504, 92.79188, 92.63555, 92.29731, 91.84467, 91.48444, 92.08432,
    91.29365, 87.45621, 84.83472, 83.09105, 81.65369, 80.13597, 79.02223,
    79.77081, 80.51665, 79.47231, 73.86306, 73.90496, 72.10558, 62.14823,
    48.79753, 45.2466,
  97.05881, 98.21315, 98.29199, 98.78909, 97.89198, 96.01106, 95.19691,
    95.94165, 96.11029, 96.48275, 96.53267, 96.66556, 95.76765, 93.41106,
    90.26992, 88.01665, 85.32555, 82.92034, 81.10154, 80.45769, 80.3614,
    78.04456, 74.85469, 69.03316, 72.25171, 77.70126, 68.54337, 49.81977,
    45.32522, 43.75951,
  97.00227, 97.86481, 99.73937, 99.8122, 101.0993, 99.72234, 98.161,
    97.30518, 96.79333, 97.14723, 96.71416, 91.70422, 90.75977, 89.36842,
    86.99384, 84.15704, 81.73763, 77.74534, 73.36809, 70.62284, 71.64487,
    67.37601, 59.71712, 55.9509, 57.21918, 56.28864, 49.66483, 45.10005,
    44.64821, 43.73959,
  98.36028, 95.48435, 98.28703, 99.63954, 98.84409, 97.31759, 96.24563,
    93.49776, 90.66312, 90.3828, 89.79199, 84.86169, 85.07793, 84.49037,
    79.93697, 76.08732, 71.48576, 68.31929, 65.67825, 64.84646, 65.92464,
    61.88798, 54.96769, 60.34003, 62.93101, 50.71669, 45.2135, 45.8013,
    45.14149, 44.18875,
  104.0159, 104.6859, 105.971, 106.3666, 104.8126, 101.6241, 94.97513,
    91.77236, 92.49879, 90.29023, 90.92115, 90.30472, 90.31901, 90.16805,
    87.55962, 78.71048, 75.58495, 71.42973, 68.47842, 69.37759, 67.23533,
    59.52382, 55.56524, 56.51432, 56.91095, 48.98024, 46.11179, 46.27785,
    46.18746, 44.78746,
  97.91975, 98.65234, 98.73934, 96.77921, 95.51065, 94.98725, 95.13709,
    95.75871, 93.38314, 93.34023, 93.72685, 91.81117, 92.84726, 93.22704,
    90.10096, 86.03109, 82.15632, 79.5621, 78.55614, 76.83794, 66.07954,
    59.14167, 58.35457, 51.40405, 47.95071, 47.09743, 45.68521, 45.06791,
    45.19296, 44.5594,
  91.63749, 92.12445, 91.84206, 91.32108, 91.27137, 92.48068, 96.15699,
    97.53819, 94.81232, 94.51504, 94.07026, 93.55514, 93.24129, 91.90634,
    89.71807, 85.82564, 82.02237, 79.61944, 79.12679, 74.52289, 60.81959,
    56.92722, 50.55656, 48.24987, 47.21947, 46.74244, 45.62201, 44.86605,
    44.43791, 44.04552,
  93.17038, 94.09597, 94.50034, 94.25423, 94.0153, 95.00394, 95.99551,
    96.14017, 95.91285, 94.55315, 93.81057, 91.95888, 90.8873, 90.93687,
    88.49303, 85.25437, 80.02042, 72.11506, 68.88271, 64.14803, 52.97952,
    51.8388, 49.08904, 48.08051, 47.44246, 46.63657, 45.57123, 44.90977,
    44.49676, 44.02987,
  92.88631, 93.24256, 93.24646, 93.36375, 93.9881, 93.79835, 94.41454,
    95.39909, 94.81067, 93.88779, 92.4814, 92.46465, 93.2821, 91.20207,
    87.25397, 80.55608, 74.06674, 68.22231, 68.5347, 65.34029, 51.87682,
    51.95064, 49.7005, 48.13499, 46.97668, 46.58529, 45.44994, 44.33628,
    44.18161, 43.96281,
  90.88212, 92.24595, 92.1281, 92.56578, 92.68598, 93.09216, 93.31645,
    93.80875, 94.23215, 93.15687, 92.98114, 93.17661, 92.26633, 90.87278,
    88.7999, 80.91368, 69.50025, 64.2803, 66.18447, 62.03894, 52.17316,
    50.95272, 49.01587, 47.575, 45.87564, 45.52231, 45.05042, 44.04143,
    43.90324, 43.7871,
  88.54554, 88.03281, 86.90153, 87.51419, 89.43356, 90.53342, 92.1898,
    92.82982, 92.60789, 92.39767, 92.74306, 92.02925, 86.19847, 87.68335,
    87.5124, 84.531, 82.55788, 80.78225, 80.26181, 73.42124, 60.22435,
    52.13107, 48.58897, 47.29124, 45.45027, 44.8797, 44.62437, 44.09175,
    43.86039, 43.77497,
  81.55737, 81.28781, 80.84987, 80.99319, 83.1255, 85.21969, 87.2744,
    88.64947, 89.66193, 92.3161, 91.39331, 84.51167, 83.19339, 82.92397,
    81.41824, 78.59863, 77.42785, 76.46476, 74.8173, 72.38999, 64.86153,
    55.94159, 49.82734, 48.01127, 46.24018, 45.07908, 44.5501, 44.12832,
    43.86708, 43.76638,
  76.48859, 76.18085, 75.30179, 75.39841, 76.86882, 78.60559, 80.31533,
    81.57737, 82.82048, 84.00053, 80.20966, 75.14935, 75.80937, 74.74496,
    72.01767, 68.33218, 66.11812, 64.8746, 64.86221, 63.5905, 61.60017,
    59.45789, 54.57249, 50.39865, 47.49334, 45.72242, 44.57815, 44.13012,
    43.8749, 43.77972,
  76.81287, 73.55767, 72.55668, 72.45029, 73.11327, 73.15382, 74.03146,
    74.35397, 76.1068, 75.46692, 70.00443, 67.27869, 67.71514, 66.5822,
    64.73298, 62.73477, 60.47995, 59.05932, 58.4817, 57.55615, 58.21364,
    59.14407, 57.94971, 56.58666, 51.63864, 46.91803, 44.83004, 44.4045,
    43.90532, 43.76528,
  76.57142, 74.79964, 72.92973, 72.50065, 74.10198, 74.51719, 73.07593,
    71.06899, 71.17102, 68.96134, 64.38639, 64.44422, 64.70528, 64.20446,
    62.61557, 61.46838, 59.75672, 56.92936, 55.5092, 54.9225, 55.50806,
    56.22244, 54.52468, 54.8259, 54.21947, 49.34728, 45.67116, 45.30085,
    44.46933, 43.83932,
  84.02925, 82.87633, 82.23975, 81.96562, 81.77481, 80.6964, 80.34402,
    79.18043, 78.32616, 72.79192, 68.26733, 69.70412, 69.86926, 69.27441,
    67.21096, 64.76817, 62.601, 59.67242, 56.51908, 55.38427, 55.51134,
    55.08538, 53.52055, 52.3918, 52.37619, 52.04771, 48.6915, 45.97874,
    45.17413, 44.20356,
  88.16456, 90.40295, 85.79375, 84.60587, 85.29226, 84.54533, 82.23651,
    81.00174, 81.7566, 77.59583, 72.10698, 73.17152, 72.83153, 71.14672,
    68.49805, 65.91193, 62.92751, 60.67448, 57.68925, 54.99545, 54.57663,
    54.17727, 52.71945, 51.31096, 50.25091, 51.11184, 51.12158, 48.47106,
    46.98165, 45.32961,
  95.73248, 99.73769, 96.83579, 93.06757, 90.85438, 88.69715, 88.31265,
    87.021, 82.46302, 77.52516, 75.08793, 74.90382, 74.03689, 70.65305,
    66.84138, 64.4426, 62.23505, 60.32514, 58.1715, 55.79998, 55.44083,
    55.12371, 52.82513, 50.9589, 50.46545, 50.61357, 51.51018, 49.79691,
    46.50879, 44.97676,
  97.25124, 99.11266, 94.33672, 92.05786, 91.09514, 88.74869, 88.29,
    85.61774, 79.8297, 76.67307, 76.28011, 75.88866, 74.29419, 71.1052,
    68.21071, 65.54319, 63.45547, 62.47552, 61.12579, 59.68351, 60.77671,
    62.46906, 61.24287, 57.54251, 54.99259, 54.08372, 54.72976, 53.3448,
    47.17955, 43.94907,
  96.09297, 97.31855, 95.28372, 95.07843, 95.13573, 92.52694, 89.52456,
    84.79538, 79.57456, 79.4379, 79.13438, 78.95187, 77.79759, 75.37821,
    73.49043, 70.93726, 68.24895, 67.20802, 66.49167, 65.97478, 65.91256,
    64.06322, 60.53928, 58.04487, 56.37472, 55.54977, 54.78121, 56.16251,
    53.18634, 45.83594,
  89.68842, 90.37514, 93.97852, 96.74339, 96.42749, 95.32592, 90.048,
    82.22832, 79.44112, 79.99371, 79.1318, 78.55471, 78.02772, 77.55253,
    76.64691, 74.19721, 71.22338, 68.66742, 64.92377, 61.02706, 59.22098,
    57.17831, 54.82459, 53.13757, 52.74254, 52.53003, 51.64552, 50.04007,
    49.53366, 46.81989,
  87.2306, 88.6123, 89.67123, 89.73494, 89.98146, 92.11813, 90.74125,
    82.79668, 78.82989, 80.5488, 81.24612, 81.08946, 79.58372, 77.44439,
    73.88902, 68.93177, 63.3349, 58.40134, 56.09484, 53.73825, 51.78002,
    51.00897, 50.23162, 49.47425, 49.07543, 49.16059, 48.59385, 46.99787,
    45.31557, 43.93211,
  44.18567, 44.29854, 44.39737, 44.50831, 44.55101, 44.66157, 44.80256,
    44.96413, 45.17411, 45.4564, 46.48579, 46.65849, 45.12902, 45.42017,
    45.65952, 45.28581, 45.2714, 45.56727, 45.92315, 46.7708, 47.31607,
    46.87716, 47.223, 48.19802, 48.84655, 48.59296, 51.25267, 52.63086,
    46.77462, 44.9204,
  45.90436, 46.16008, 45.94139, 46.39693, 46.27977, 46.2281, 46.52509,
    46.76575, 47.01112, 47.33574, 47.78651, 48.48681, 49.05206, 48.23267,
    47.70509, 48.07795, 47.65155, 48.13733, 48.98977, 49.80005, 50.00161,
    49.98341, 50.51801, 51.94249, 56.5592, 57.55172, 51.50106, 53.93554,
    47.56802, 45.66522,
  47.21722, 47.41816, 47.58042, 47.84504, 48.02728, 48.23339, 48.4824,
    48.77652, 49.08876, 49.40531, 49.77163, 50.4131, 51.00309, 51.89991,
    52.48369, 51.77638, 52.05381, 52.94681, 53.4946, 54.34584, 55.95061,
    57.78959, 58.56803, 57.82475, 61.16885, 63.14245, 54.85175, 53.12302,
    47.58263, 46.37215,
  50.53063, 51.03599, 51.6229, 52.27277, 52.90203, 53.77067, 54.0464,
    53.87056, 54.18828, 54.63443, 54.89648, 55.56539, 55.75928, 55.4536,
    56.94238, 58.31367, 57.49302, 56.21511, 57.02729, 58.04276, 60.43013,
    60.96556, 58.71644, 63.22841, 65.11366, 58.25356, 57.55281, 52.26461,
    47.68957, 45.43842,
  55.23945, 55.37172, 56.00871, 56.65401, 57.03162, 57.30312, 57.45851,
    57.46308, 58.12299, 58.62712, 58.36253, 58.70026, 58.97316, 59.44071,
    59.80105, 60.23748, 59.44341, 57.7321, 57.87555, 62.87851, 64.7933,
    56.23911, 56.28717, 57.66314, 59.45107, 58.54096, 54.90051, 55.28107,
    54.64672, 47.87436,
  58.68223, 59.50533, 60.5966, 62.02061, 61.93364, 61.53613, 62.3232,
    62.69694, 62.60133, 63.21692, 64.11686, 66.61233, 69.32201, 68.58201,
    67.6177, 76.3904, 86.45473, 71.37781, 60.66895, 61.21212, 58.35675,
    54.63509, 55.51624, 56.84879, 59.23337, 58.02631, 61.29388, 77.67965,
    68.92628, 46.59003,
  63.56348, 65.1292, 66.70194, 68.41622, 68.94427, 69.41437, 71.07124,
    72.85533, 72.33247, 71.15587, 70.45419, 68.37216, 65.31129, 64.83138,
    69.00021, 74.88001, 69.8923, 62.04022, 58.25532, 57.71341, 55.89644,
    54.83721, 55.59144, 58.02198, 58.93383, 55.19923, 64.2754, 81.24816,
    65.34341, 44.6308,
  68.50381, 70.14082, 71.47421, 72.64538, 71.95556, 72.84721, 73.81519,
    69.07647, 65.04906, 63.88189, 62.19338, 60.32811, 58.8194, 58.66011,
    59.22766, 59.91825, 59.80001, 58.72226, 55.83641, 55.18852, 54.34343,
    54.25836, 55.93203, 57.89585, 56.71318, 54.37935, 65.00137, 70.20221,
    51.50658, 45.3393,
  71.49285, 71.64331, 71.83033, 70.90388, 69.14702, 68.74846, 65.44701,
    63.0624, 62.99225, 62.51712, 61.77542, 61.0407, 60.81099, 64.60284,
    67.14764, 61.88349, 60.8327, 62.09916, 61.6055, 58.45498, 56.17339,
    58.62481, 63.17187, 62.93089, 57.61367, 58.02456, 60.61567, 56.9242,
    47.39864, 45.05927,
  78.4574, 79.82532, 79.50635, 79.45839, 76.73029, 70.81007, 64.90945,
    66.24614, 66.82117, 68.56461, 70.52343, 73.69695, 73.57561, 70.48222,
    66.70477, 67.74116, 68.33106, 67.56154, 65.11723, 63.44944, 63.81558,
    62.99476, 61.77457, 57.8207, 65.36124, 79.19524, 64.8818, 48.04265,
    45.23097, 44.0075,
  84.90586, 83.5932, 83.0097, 81.86232, 81.33319, 80.91657, 80.35748,
    80.55421, 81.05873, 82.51762, 83.743, 71.09846, 66.86409, 66.0396,
    65.59661, 65.60452, 65.7846, 64.71846, 62.79211, 61.47739, 62.8881,
    60.70324, 55.33134, 51.98165, 53.76552, 55.06623, 49.3518, 44.85975,
    44.52137, 43.93448,
  91.85854, 86.40234, 89.09131, 88.81401, 87.50119, 85.58971, 84.31917,
    81.50058, 78.82288, 79.1392, 76.27562, 67.93525, 69.33424, 68.54039,
    63.89061, 63.35173, 61.07156, 59.67901, 58.02999, 57.29011, 58.56797,
    56.41936, 50.59069, 55.17072, 58.23778, 47.87852, 44.69634, 45.09717,
    44.81253, 44.21201,
  99.31786, 98.08864, 99.77988, 97.96094, 95.15037, 90.28105, 82.54266,
    78.70408, 79.09192, 77.41795, 77.83183, 73.0301, 74.77026, 75.23821,
    66.31396, 61.5496, 59.87068, 58.14326, 56.45391, 57.63963, 57.82428,
    53.55651, 50.19508, 53.57703, 55.61153, 46.82806, 45.25844, 45.39563,
    45.40325, 44.59676,
  95.80243, 97.78989, 95.11353, 90.69469, 86.97533, 84.84525, 83.91326,
    83.24635, 80.72068, 79.6472, 80.67011, 79.7579, 81.61385, 84.43378,
    87.56542, 72.08466, 61.08913, 62.11561, 62.19696, 61.15576, 56.29149,
    54.68668, 57.29659, 50.21155, 47.08662, 46.13989, 45.22581, 44.79155,
    44.89392, 44.47738,
  86.33148, 84.66566, 82.84103, 80.82198, 79.439, 81.00105, 85.77277,
    84.89729, 81.54972, 80.75269, 79.90095, 79.48849, 78.56491, 81.79292,
    82.83893, 66.85131, 65.2062, 62.71015, 63.24402, 64.295, 60.31303,
    53.8429, 48.37693, 46.57037, 46.01474, 46.03733, 45.22707, 44.65416,
    44.38748, 44.14059,
  82.71271, 81.521, 81.01714, 80.02229, 79.27904, 79.61252, 80.22347,
    79.82719, 79.05173, 78.14297, 78.11642, 73.72153, 69.61086, 70.06413,
    66.6173, 63.51133, 62.18167, 58.76662, 57.80106, 56.14919, 49.90901,
    48.38274, 46.47372, 46.04702, 46.11909, 45.90997, 45.23604, 44.69876,
    44.40631, 44.11819,
  81.52176, 80.34928, 79.61369, 78.85979, 78.65177, 77.9035, 77.9418,
    78.63215, 77.55032, 75.20535, 70.35222, 69.66353, 71.88155, 66.7932,
    63.06388, 60.6134, 58.06452, 55.57757, 56.50038, 55.34388, 47.62917,
    48.0825, 47.04501, 46.16195, 45.83554, 45.89248, 45.17683, 44.386,
    44.21995, 44.07721,
  77.5378, 76.83569, 75.05322, 74.26267, 73.11129, 72.80575, 72.22457,
    71.59788, 71.2459, 68.38895, 68.49574, 70.02964, 67.61392, 65.58644,
    65.45714, 60.74421, 55.10144, 52.54665, 54.8147, 53.67404, 48.02668,
    47.96541, 47.10667, 46.27687, 45.34803, 45.23843, 44.87666, 44.17418,
    44.06514, 43.97425,
  75.02467, 73.07732, 69.76893, 67.62472, 66.99915, 66.04754, 65.57639,
    65.45644, 64.35318, 63.50339, 64.96439, 63.43874, 58.56014, 58.9672,
    59.20574, 58.38285, 58.80304, 59.69831, 61.92462, 60.65679, 54.08549,
    49.23473, 46.77872, 46.24783, 45.09574, 44.74319, 44.5715, 44.18357,
    44.03671, 43.96422,
  70.74303, 68.64882, 65.70499, 63.09769, 62.3833, 61.79405, 61.33435,
    60.93015, 60.73029, 62.5088, 62.77201, 58.45457, 57.43208, 57.84257,
    57.80153, 57.25911, 58.19911, 59.57181, 60.12566, 59.91297, 56.24372,
    51.03441, 47.22718, 46.53772, 45.53917, 44.81344, 44.50259, 44.22063,
    44.04401, 43.96826,
  67.35322, 65.54331, 62.72743, 60.53094, 59.70064, 59.29686, 59.0327,
    58.96585, 59.69706, 61.40592, 59.82, 56.7041, 57.80247, 57.99206,
    57.01683, 55.38685, 54.65478, 54.07777, 54.10077, 53.50671, 52.33787,
    51.54001, 49.56211, 47.65482, 46.2172, 45.25915, 44.52343, 44.22032,
    44.06172, 43.97346,
  67.32045, 64.15614, 61.86766, 60.31707, 59.62214, 58.6659, 58.56169,
    58.35929, 59.84381, 60.43697, 57.07012, 54.93275, 55.35275, 54.74562,
    53.65469, 52.60285, 51.38154, 50.51826, 50.23627, 49.66737, 50.91329,
    52.01664, 50.41322, 50.91476, 48.62187, 45.98212, 44.67637, 44.37923,
    44.08127, 43.97476,
  66.0177, 64.31718, 61.93049, 60.43317, 60.77184, 60.68459, 59.56808,
    57.96221, 58.08186, 56.73791, 53.08443, 52.43566, 52.43412, 52.19174,
    51.36649, 51.21345, 50.86498, 49.51763, 48.83799, 48.50594, 49.53656,
    50.3032, 48.37629, 49.46987, 49.78304, 47.24088, 45.01583, 44.86931,
    44.40712, 44.02313,
  66.25344, 65.12181, 63.95286, 63.09414, 62.37481, 61.12102, 60.61453,
    59.8245, 59.63158, 56.01617, 52.0819, 52.55249, 52.92865, 53.20723,
    52.75413, 52.29075, 52.00587, 50.87013, 49.18037, 48.53567, 48.51023,
    48.39844, 47.80573, 47.65445, 48.28384, 48.52064, 46.72342, 45.21299,
    44.80451, 44.24154,
  66.0273, 66.19518, 63.04015, 61.51157, 61.34624, 60.50697, 59.06891,
    58.52778, 59.68481, 56.96813, 52.57084, 53.33799, 53.87393, 53.9054,
    53.44379, 53.03057, 52.17253, 51.61652, 50.29328, 48.72508, 48.54422,
    48.60394, 48.20257, 47.42422, 46.81363, 47.7823, 47.99105, 46.53146,
    45.89017, 44.93755,
  67.24804, 68.54305, 66.66991, 63.8837, 62.03462, 60.58162, 60.98126,
    61.55132, 59.51884, 56.10706, 54.298, 54.76095, 55.24059, 54.31958,
    52.92966, 52.43665, 51.9388, 51.45852, 50.56469, 49.14348, 48.96748,
    49.03786, 47.92944, 47.01642, 46.99086, 47.36207, 48.31124, 47.58131,
    45.7108, 44.71018,
  68.33788, 68.71771, 65.40808, 63.04655, 61.92603, 60.27889, 60.97682,
    60.66648, 57.28141, 54.78934, 54.65248, 54.9072, 54.76022, 53.69868,
    52.80326, 52.02397, 51.26476, 51.085, 50.52758, 49.46532, 49.96876,
    51.50146, 51.71361, 50.20369, 49.27268, 49.12415, 50.11465, 49.80891,
    46.04495, 44.02302,
  68.02382, 67.19701, 64.78086, 63.68673, 63.21905, 61.831, 61.05344,
    58.77494, 54.96116, 54.24121, 53.86992, 53.9319, 53.85179, 53.30428,
    53.30417, 52.87137, 52.02623, 52.07851, 52.39546, 52.63187, 53.24395,
    53.19938, 51.84547, 50.6527, 50.00904, 49.92294, 49.85257, 51.36993,
    49.81145, 45.21644,
  65.52669, 63.97216, 64.09906, 64.49633, 64.04171, 64.0508, 61.53654,
    56.56455, 53.91347, 53.75826, 52.92544, 52.80108, 53.18303, 53.93099,
    55.04313, 55.54935, 55.45352, 55.33715, 54.06715, 52.28928, 51.66303,
    50.82243, 49.61953, 48.78814, 48.7397, 48.882, 48.66967, 47.99177,
    47.96329, 46.03112,
  64.73904, 64.19382, 63.54854, 62.36726, 61.94352, 63.7711, 63.92814,
    58.83738, 55.65017, 56.47813, 57.17915, 57.90452, 58.13667, 58.03885,
    57.5766, 56.58507, 54.62486, 52.42272, 51.30785, 49.85012, 48.72713,
    48.30228, 47.8776, 47.4435, 47.18991, 47.35823, 47.05004, 46.14825,
    45.23106, 44.19022,
  31.21135, 31.26128, 31.30381, 31.3622, 31.36663, 31.39029, 31.42309,
    31.47893, 31.61026, 31.77498, 32.65834, 32.77625, 31.60489, 31.7891,
    31.93258, 31.58587, 31.47986, 31.5797, 31.70495, 32.30421, 32.63241,
    32.17508, 32.28576, 32.97128, 33.44476, 33.26427, 35.7197, 37.07351,
    33.14369, 31.86181,
  32.0137, 32.12721, 31.92243, 32.23438, 32.07856, 31.94452, 32.08078,
    32.18184, 32.30536, 32.4942, 32.8288, 33.32064, 33.62715, 32.9175,
    32.50136, 32.64038, 32.17974, 32.38876, 32.98219, 33.51436, 33.59363,
    33.39647, 33.80144, 34.81161, 39.21036, 40.47346, 35.93261, 38.20842,
    33.74387, 32.31145,
  32.6692, 32.7461, 32.74836, 32.83332, 32.85909, 32.87471, 32.91561,
    33.02339, 33.12699, 33.19557, 33.26991, 33.56744, 33.78996, 34.22468,
    34.46908, 33.82738, 33.91194, 34.52019, 34.83152, 35.39827, 36.62986,
    38.13347, 39.16687, 38.72152, 43.1344, 45.80486, 38.09141, 37.66268,
    33.71261, 32.83509,
  34.74739, 34.95292, 35.25162, 35.58039, 35.94108, 36.53695, 36.63267,
    36.28998, 36.29628, 36.42595, 36.32373, 36.41172, 36.05138, 35.51619,
    36.57117, 37.73504, 37.25441, 36.40082, 37.07833, 37.94457, 40.21645,
    41.23581, 39.69753, 44.64943, 46.93957, 40.71291, 40.40067, 36.94722,
    33.69633, 32.21893,
  38.79986, 38.89825, 39.31243, 39.77558, 40.05974, 40.2492, 40.30251,
    40.18154, 40.5318, 40.56293, 39.79398, 39.17661, 38.53342, 38.43038,
    38.83309, 39.39382, 38.87914, 38.2333, 38.62697, 43.55956, 45.3235,
    38.47071, 38.40876, 39.85747, 41.40608, 40.32275, 37.91548, 37.99441,
    38.06129, 33.89417,
  42.90058, 43.57038, 44.39814, 45.41026, 45.15688, 44.71535, 45.19844,
    45.29093, 44.93603, 44.78579, 44.33955, 45.05049, 45.9599, 45.01274,
    43.71685, 52.32983, 62.2427, 49.8904, 41.43474, 42.59351, 40.41782,
    37.04313, 37.54607, 38.30645, 40.39988, 39.45823, 43.16539, 57.80903,
    50.71184, 32.98863,
  47.02876, 48.1286, 49.18805, 50.40186, 50.6656, 51.01481, 52.68718,
    54.56059, 54.46204, 53.56127, 52.64023, 50.03045, 46.55185, 45.05482,
    49.70477, 56.84912, 52.01648, 43.36544, 40.18821, 39.5807, 37.96053,
    37.05503, 37.59616, 39.55823, 40.74783, 37.73632, 48.07997, 65.44596,
    49.62307, 31.52893,
  51.37611, 53.00611, 54.46518, 56.05602, 56.31071, 58.11394, 60.13454,
    57.46689, 54.6095, 53.14012, 50.66042, 47.15626, 43.75416, 41.98149,
    42.20517, 42.76093, 41.74195, 40.4124, 38.26505, 37.76216, 37.06791,
    36.83831, 38.1291, 39.88768, 39.35044, 37.16198, 48.85681, 54.63733,
    37.41284, 32.54436,
  57.28215, 58.49558, 59.37911, 59.51868, 59.15963, 59.5674, 57.29989,
    55.01052, 53.99476, 52.21817, 49.53976, 46.31129, 43.49374, 44.77083,
    45.68686, 41.43769, 40.85231, 42.07626, 41.80735, 39.37539, 37.60493,
    39.36913, 43.15866, 43.14913, 39.43686, 39.56316, 45.21817, 44.38139,
    34.54964, 32.41622,
  62.70608, 64.76356, 65.06557, 65.43553, 63.84621, 59.18777, 54.08834,
    53.87799, 53.08382, 52.36076, 51.93561, 52.82884, 51.01286, 47.50609,
    44.01593, 44.01634, 44.66953, 44.46022, 43.06392, 42.74908, 43.2991,
    43.594, 43.59865, 41.04824, 48.51636, 59.9284, 48.87125, 35.67612,
    32.68859, 31.34707,
  86.04472, 88.80721, 80.85294, 70.79814, 68.69854, 65.08864, 60.99316,
    62.541, 63.34598, 71.93574, 77.40908, 53.087, 45.40683, 43.30595,
    42.28959, 43.10484, 43.88056, 43.63661, 42.41751, 42.09733, 44.59621,
    43.65374, 39.54141, 36.95375, 40.15923, 42.93, 36.97012, 32.14667,
    31.7833, 31.21622,
  96.76215, 92.74481, 95.72607, 96.93104, 94.46577, 80.76964, 80.16541,
    72.82803, 62.01843, 64.2823, 61.60743, 46.94237, 47.05408, 46.58442,
    42.4092, 42.61417, 41.38445, 40.93151, 39.98394, 40.00185, 42.52975,
    40.95749, 35.92469, 40.26144, 42.44215, 34.4373, 31.80456, 32.22904,
    32.05263, 31.46753,
  100.1492, 101.1091, 105.1807, 106.5369, 106.3127, 103.4259, 88.85235,
    65.71688, 64.57746, 59.046, 56.2485, 47.95767, 50.33299, 51.65811,
    44.39416, 42.34357, 41.60545, 40.3129, 39.13132, 41.09222, 42.25834,
    38.50448, 35.43663, 40.06309, 41.57404, 33.58646, 32.18644, 32.42722,
    32.62543, 31.80298,
  101.7161, 106.7374, 106.7372, 104.3947, 101.7179, 98.34703, 94.80344,
    95.06518, 84.67464, 80.38145, 86.97507, 79.68937, 78.00829, 74.37238,
    63.258, 50.15246, 41.78896, 43.28268, 44.36341, 44.81693, 41.03531,
    39.99215, 42.176, 36.90668, 34.16803, 32.95402, 32.19096, 31.87236,
    32.18081, 31.72863,
  89.49129, 89.52451, 83.81065, 79.41049, 75.10043, 86.14627, 96.93047,
    97.55764, 95.17135, 94.91097, 86.7042, 67.22723, 52.98945, 57.57751,
    61.51794, 46.13483, 45.79357, 45.23102, 48.3454, 49.65294, 44.36769,
    39.78238, 35.73416, 33.50806, 32.74362, 32.99652, 32.25664, 31.76387,
    31.64687, 31.40358,
  72.71319, 70.75528, 69.70433, 68.69706, 69.23254, 73.57436, 77.76678,
    74.76159, 70.5892, 65.30826, 59.48203, 52.33395, 46.3676, 48.37423,
    47.24523, 45.00791, 45.60029, 43.40453, 44.10109, 43.36585, 37.11773,
    34.81935, 33.0009, 32.79085, 33.05412, 32.8719, 32.29658, 31.83238,
    31.61377, 31.34638,
  68.06772, 66.67277, 65.77576, 65.56189, 65.87229, 65.10004, 64.28304,
    63.4192, 60.46471, 56.3419, 50.44234, 49.15552, 51.34273, 47.60258,
    44.70932, 43.98812, 42.64632, 40.57488, 42.71854, 41.56821, 33.8191,
    34.16574, 33.612, 32.9479, 32.75407, 32.85964, 32.21584, 31.55045,
    31.44877, 31.31383,
  63.95418, 63.84851, 62.61434, 62.05413, 60.99147, 60.35381, 59.66439,
    59.15012, 57.44223, 52.66803, 50.52076, 51.11666, 48.78827, 47.16441,
    48.34795, 45.16868, 40.01218, 37.50687, 40.85411, 39.94184, 34.25906,
    34.41153, 33.92355, 33.2159, 32.29668, 32.33288, 31.9993, 31.36216,
    31.27906, 31.22608,
  63.22479, 62.27501, 59.72658, 58.00062, 57.34193, 56.48726, 55.89586,
    55.42136, 53.21296, 50.21478, 49.9124, 47.13224, 41.23826, 41.16133,
    41.67572, 40.80667, 40.97947, 41.83653, 45.04987, 44.34016, 38.45692,
    35.29812, 33.91108, 33.24957, 32.14575, 31.91532, 31.75894, 31.37761,
    31.26638, 31.21809,
  60.85851, 59.88989, 57.72255, 55.44134, 54.88707, 54.36533, 53.78482,
    52.68964, 50.80252, 50.38297, 48.21623, 41.60907, 38.47776, 38.30994,
    38.1944, 37.69852, 39.20417, 41.42048, 43.56825, 44.56282, 41.5421,
    37.30567, 34.36275, 33.45928, 32.55766, 31.97393, 31.69459, 31.42425,
    31.28854, 31.2231,
  58.43968, 58.22576, 55.80779, 53.88779, 53.17081, 52.67819, 51.94275,
    50.70158, 49.44215, 48.74266, 44.03498, 38.28802, 38.13099, 38.45962,
    38.08787, 37.19726, 37.24526, 37.58825, 38.76836, 39.23623, 38.70103,
    38.14254, 36.41953, 34.37317, 33.04621, 32.3032, 31.70681, 31.42006,
    31.32043, 31.24997,
  58.56114, 56.44339, 54.36914, 53.04097, 52.24564, 51.20976, 50.63604,
    49.4477, 49.30663, 47.41294, 41.31834, 37.57293, 37.66797, 37.53362,
    37.08113, 36.52, 35.80342, 35.47579, 35.55463, 35.24873, 36.64546,
    37.54947, 37.16055, 37.71925, 35.57481, 33.04985, 31.87119, 31.59764,
    31.33844, 31.25672,
  56.63459, 55.42986, 53.16282, 51.84512, 52.28123, 52.57719, 51.86079,
    50.10631, 49.3862, 45.73599, 39.4493, 37.17428, 36.7527, 36.50632,
    35.90675, 36.05306, 35.8618, 34.76816, 34.25315, 34.10138, 35.48426,
    35.99466, 34.81035, 36.45328, 36.93943, 34.27097, 32.15219, 32.07266,
    31.65791, 31.28512,
  55.67796, 54.95037, 54.0577, 53.68987, 53.65902, 53.50218, 53.75826,
    53.20591, 52.1839, 45.94365, 38.96691, 37.50272, 37.14387, 37.27262,
    36.9993, 36.87792, 37.03839, 36.11027, 34.56102, 34.23556, 34.64838,
    34.64267, 34.12773, 34.31356, 35.4693, 35.72812, 33.84846, 32.45975,
    32.06305, 31.47502,
  55.92146, 56.97372, 54.19404, 53.2469, 53.69635, 53.67297, 52.92002,
    52.3411, 52.25233, 46.31932, 38.88142, 37.67233, 37.63965, 37.64643,
    37.53192, 37.56181, 37.21913, 37.05776, 35.68841, 34.2029, 34.45936,
    34.81991, 34.68533, 33.86045, 33.26889, 34.53795, 34.8295, 33.48661,
    33.08494, 32.06078,
  57.06163, 59.09419, 57.66078, 55.56815, 54.00986, 52.97866, 53.87471,
    54.37453, 51.01044, 44.7148, 39.71021, 38.53362, 38.76104, 38.00343,
    37.04493, 36.96335, 36.84346, 36.9253, 36.07755, 34.63263, 34.99063,
    35.41399, 34.31921, 33.28392, 33.12069, 33.67676, 35.00848, 34.31464,
    32.93539, 31.91637,
  58.09569, 59.38708, 56.46804, 54.45842, 53.45613, 52.34531, 53.70699,
    53.60845, 48.58609, 43.13401, 40.15327, 38.9353, 38.42992, 37.52822,
    36.99219, 36.61891, 36.25953, 36.53716, 35.92175, 34.56212, 35.42544,
    37.40976, 37.64845, 35.93037, 34.99945, 35.04534, 36.65083, 36.58546,
    33.11501, 31.25051,
  57.52391, 57.57401, 55.40085, 54.5879, 54.73955, 54.08545, 54.25863,
    51.89472, 46.21853, 42.65474, 39.74642, 38.33374, 37.69036, 37.04895,
    37.22616, 37.01064, 36.31216, 36.41747, 36.58271, 36.51138, 38.0125,
    38.76781, 37.63708, 36.21259, 35.46672, 35.5562, 35.83485, 37.87662,
    36.37653, 32.22828,
  55.01461, 54.15842, 54.5876, 55.728, 56.45027, 57.51906, 55.7089, 50.40936,
    45.84802, 42.68587, 38.8844, 36.54901, 35.79017, 36.29683, 37.63318,
    38.38501, 38.5534, 38.93993, 37.85841, 36.31605, 36.2876, 35.84192,
    34.77709, 34.0881, 34.18745, 34.60406, 34.65654, 34.45655, 35.00562,
    32.94997,
  53.46158, 53.53756, 53.35491, 52.87127, 53.11179, 55.94889, 56.43576,
    50.50382, 45.33121, 42.98866, 40.75961, 39.52275, 39.12453, 39.74401,
    40.30199, 40.04945, 38.72504, 37.10527, 36.11869, 34.7646, 33.94906,
    33.67991, 33.44026, 33.20447, 33.17636, 33.63909, 33.68027, 33.03137,
    32.36821, 31.48538,
  31.41252, 31.46955, 31.49963, 31.53003, 31.53205, 31.52726, 31.54217,
    31.58476, 31.67506, 31.80536, 32.79342, 32.90239, 31.75217, 31.96879,
    32.11943, 31.73141, 31.58411, 31.63934, 31.72813, 32.36559, 32.68122,
    32.12987, 32.12052, 32.7661, 33.12569, 32.74058, 35.47042, 37.25195,
    33.62823, 32.25118,
  31.86638, 31.93911, 31.721, 32.03023, 31.85303, 31.67992, 31.76275,
    31.84919, 31.97054, 32.16982, 32.59097, 33.1835, 33.50525, 32.79121,
    32.45045, 32.48887, 31.92691, 32.01481, 32.58499, 33.15451, 33.13107,
    32.62748, 32.74018, 33.75631, 38.07284, 38.73828, 35.81148, 39.06515,
    34.45575, 32.84657,
  31.80177, 31.84221, 31.82227, 31.89351, 31.87299, 31.86183, 31.89826,
    31.97831, 32.08513, 32.16067, 32.29577, 32.72724, 33.06064, 33.57404,
    33.71877, 32.92604, 32.84079, 33.30465, 33.48803, 33.84834, 34.88108,
    36.38021, 37.42197, 37.01488, 41.45349, 43.78821, 38.18972, 38.49588,
    34.34968, 33.45453,
  31.92943, 31.98294, 32.22617, 32.46614, 32.78315, 33.38764, 33.47604,
    33.16037, 33.21157, 33.40647, 33.49257, 34.01735, 33.9233, 33.4549,
    34.5613, 35.62631, 34.94676, 34.01248, 34.43291, 35.1251, 37.74567,
    39.05733, 37.90254, 42.31125, 43.89786, 40.07665, 40.8, 37.81671,
    34.33073, 32.72856,
  32.66642, 32.49052, 32.84326, 33.25941, 33.57536, 33.83628, 33.8927,
    33.70271, 34.18671, 34.51202, 34.34865, 34.53574, 34.58672, 34.9894,
    35.72196, 36.36409, 35.66596, 34.91621, 35.55441, 40.37897, 41.92506,
    36.54301, 36.36995, 38.18901, 40.07, 39.5879, 37.84427, 38.45649,
    39.16247, 34.47578,
  32.94669, 33.17435, 34.01919, 35.11108, 34.91988, 34.45353, 34.78656,
    34.66489, 34.29091, 34.48852, 34.81734, 37.04423, 39.66017, 39.74519,
    39.2573, 46.57125, 53.58584, 44.53928, 38.54233, 40.32322, 38.39807,
    34.95086, 35.45577, 36.46878, 39.26909, 38.79146, 41.42303, 54.42943,
    49.9274, 33.86761,
  33.40923, 33.87736, 34.81859, 35.85808, 35.96045, 35.93158, 37.29353,
    39.18641, 39.51878, 39.76999, 40.76702, 40.43212, 39.22698, 39.49376,
    44.5648, 51.36488, 48.37154, 40.65217, 37.79206, 37.41636, 35.83361,
    34.86305, 35.52055, 38.17472, 39.78699, 37.20959, 46.90069, 62.26871,
    49.14259, 32.30513,
  34.10607, 34.8096, 36.09993, 37.46035, 37.62326, 39.96348, 42.71515,
    40.71305, 39.07032, 39.36371, 39.38798, 38.33241, 37.15917, 37.2973,
    39.07831, 40.39323, 39.41267, 38.0039, 36.07178, 35.66675, 35.03651,
    34.83961, 36.42048, 39.0617, 38.60583, 36.8409, 49.18007, 54.36728,
    38.64529, 32.59084,
  36.96578, 37.59975, 38.97907, 39.56171, 40.06668, 41.85106, 40.83035,
    39.24244, 39.28506, 39.28135, 38.66031, 37.55947, 36.81978, 40.34161,
    42.4798, 38.61699, 38.1866, 39.67058, 39.65843, 37.26136, 35.25513,
    37.08158, 41.79934, 42.36025, 38.4496, 39.18373, 45.46333, 43.52362,
    34.71043, 32.52362,
  41.51422, 43.58982, 45.42965, 47.2044, 46.72301, 42.43938, 37.96053,
    38.00068, 37.77573, 37.74352, 39.22169, 43.09337, 44.44776, 43.19732,
    40.95126, 40.98816, 41.83211, 42.29671, 40.63077, 39.1651, 39.494,
    40.2014, 41.08328, 39.10753, 45.11982, 55.51937, 47.39198, 35.80972,
    33.00156, 31.68968,
  55.89689, 58.44576, 54.17729, 48.45197, 47.00118, 44.94873, 41.32525,
    43.34546, 45.47102, 53.81099, 58.24356, 43.4857, 39.56281, 39.00413,
    38.38154, 39.09435, 40.17072, 40.15404, 39.16162, 39.21148, 41.86182,
    41.39704, 37.92658, 35.72813, 39.69255, 43.34319, 37.47294, 32.5594,
    32.12569, 31.53864,
  70.09546, 58.52769, 61.62629, 63.88789, 61.33881, 53.09554, 55.2051,
    51.64217, 45.35822, 49.52015, 49.1628, 37.86327, 39.25414, 40.20609,
    38.29852, 38.67093, 38.04303, 38.0197, 37.34386, 37.91706, 41.02718,
    39.81174, 35.3379, 39.06544, 40.88549, 34.4768, 32.11416, 32.53738,
    32.39119, 31.75608,
  82.72105, 80.78213, 98.87999, 102.4082, 98.10238, 84.99236, 65.74177,
    47.17777, 46.35042, 43.64202, 41.71672, 37.47422, 42.09693, 44.4242,
    39.94788, 38.96161, 38.9884, 37.89732, 36.96888, 39.25963, 40.90429,
    37.69612, 34.86119, 39.75452, 40.88229, 33.73246, 32.37481, 32.68835,
    32.93752, 32.05262,
  90.38415, 109.2217, 110.6207, 105.2391, 90.10088, 77.80119, 70.65182,
    67.20332, 56.96955, 52.94041, 60.95278, 59.90412, 62.76102, 62.36201,
    55.76287, 46.01701, 39.32608, 40.67056, 42.03157, 43.06145, 40.10038,
    38.91081, 40.45296, 36.96853, 34.54269, 33.04783, 32.37574, 32.15527,
    32.55427, 31.98825,
  66.78455, 72.05553, 67.43833, 62.84813, 56.43639, 61.80069, 82.18446,
    80.37238, 70.13571, 70.59137, 68.36681, 56.52965, 48.12868, 53.59817,
    56.11687, 43.51596, 42.79491, 43.01446, 46.90059, 47.62692, 42.4455,
    39.19212, 35.92434, 33.5099, 32.81625, 33.23518, 32.49875, 32.03443,
    32.01092, 31.70457,
  51.9077, 49.68568, 48.03596, 46.20362, 46.26603, 51.55554, 58.1395,
    56.65842, 53.91622, 52.33688, 50.00333, 44.32645, 40.72623, 44.35825,
    44.43281, 42.18981, 43.47098, 42.22429, 44.05344, 43.35206, 37.21754,
    34.78758, 32.74325, 32.55299, 33.14084, 33.15995, 32.63625, 32.11124,
    31.92517, 31.641,
  46.94086, 44.42204, 43.29732, 43.24261, 44.45417, 45.29685, 45.78689,
    46.14898, 45.41449, 44.26785, 41.11289, 41.63124, 46.0994, 44.01884,
    42.06651, 41.95943, 41.41359, 39.96629, 42.47979, 40.89437, 33.78023,
    33.9732, 33.40618, 32.72084, 32.79044, 33.09345, 32.52676, 31.8589,
    31.78791, 31.62026,
  42.5523, 41.96252, 41.64255, 42.20338, 42.33569, 42.67756, 42.60295,
    42.55091, 42.52006, 40.52465, 41.1756, 44.83073, 45.15809, 44.71955,
    46.18461, 43.61724, 39.18109, 37.17759, 40.78319, 39.41261, 34.04777,
    34.33618, 33.8793, 33.1142, 32.43345, 32.6314, 32.25229, 31.66775,
    31.61304, 31.52755,
  43.24551, 43.02604, 41.5221, 40.57598, 40.3614, 39.815, 39.51307, 39.57477,
    39.09075, 38.89928, 42.32841, 42.89251, 39.10332, 39.92373, 40.67838,
    39.68521, 39.63136, 40.64935, 43.91161, 42.63239, 37.38554, 35.105,
    34.02831, 33.35361, 32.39408, 32.21416, 32.03603, 31.64931, 31.56647,
    31.51279,
  43.69045, 42.89314, 40.81753, 38.90193, 38.46499, 38.07518, 37.88443,
    37.8171, 37.94877, 40.63697, 42.15015, 38.5699, 36.6632, 36.89893,
    36.58337, 35.96131, 37.69132, 40.35239, 42.94079, 43.68372, 40.69172,
    36.98132, 34.45677, 33.61324, 32.80516, 32.24147, 31.98033, 31.70728,
    31.57472, 31.50311,
  42.45912, 41.58164, 39.50699, 37.78341, 37.25716, 37.12475, 37.01936,
    36.96392, 37.8301, 40.31031, 38.84537, 35.37356, 36.00784, 36.57589,
    36.19518, 35.45348, 35.84903, 36.76427, 38.53519, 39.23528, 38.71161,
    38.082, 36.42217, 34.42649, 33.21036, 32.51496, 31.97502, 31.70827,
    31.61346, 31.51869,
  42.27624, 40.24956, 38.63605, 37.652, 37.09057, 36.41216, 36.29646,
    36.17855, 37.98874, 39.08108, 36.09973, 34.38693, 35.48668, 35.86513,
    35.69835, 35.37244, 34.9931, 35.01479, 35.37283, 35.30037, 36.54206,
    37.22024, 37.15667, 37.34436, 35.41834, 33.12539, 32.09749, 31.85673,
    31.66516, 31.55104,
  41.32002, 40.09584, 38.09875, 36.92678, 37.35811, 37.62353, 37.15699,
    36.41094, 37.84877, 37.42226, 34.50793, 34.30595, 35.08979, 35.34292,
    35.01838, 35.38026, 35.23857, 34.33533, 34.0008, 33.98144, 35.15908,
    35.40418, 34.96445, 36.66502, 36.92402, 34.1656, 32.34644, 32.34851,
    31.98432, 31.5824,
  40.43752, 39.50882, 38.61003, 38.22032, 38.16219, 38.14416, 38.60228,
    38.93758, 40.16166, 37.6446, 34.43311, 35.09721, 35.85342, 36.34556,
    36.2514, 36.36045, 36.46851, 35.43133, 34.19072, 34.08479, 34.32241,
    34.22323, 34.03466, 34.49045, 35.77597, 35.71019, 33.87025, 32.68836,
    32.34827, 31.72681,
  40.37164, 40.8424, 38.3389, 37.55324, 38.03775, 38.09829, 37.90532,
    38.55709, 40.82099, 38.27514, 34.67536, 35.5612, 36.45758, 36.77198,
    36.8554, 36.99618, 36.70846, 36.41928, 35.08332, 33.92862, 34.21228,
    34.38853, 34.24048, 33.60641, 33.39267, 34.73132, 34.8141, 33.50821,
    33.26385, 32.15622,
  40.86703, 42.75608, 41.4816, 39.65797, 38.27251, 37.43481, 38.75957,
    40.51081, 39.9273, 37.1106, 35.41349, 36.29864, 37.32452, 36.92072,
    36.30877, 36.33912, 36.20979, 36.28647, 35.47458, 34.27151, 34.72715,
    34.98686, 33.86605, 33.05255, 33.06972, 33.68634, 34.99675, 34.20818,
    33.08825, 31.9662,
  41.8193, 43.3848, 40.82244, 38.92402, 37.98256, 37.03209, 38.7945,
    40.09313, 37.68973, 35.62566, 35.78226, 36.65642, 37.0798, 36.5343,
    36.15138, 35.88515, 35.65849, 35.95371, 35.32544, 34.17901, 35.07349,
    36.69699, 36.63906, 35.20335, 34.68976, 34.79747, 36.4412, 36.20721,
    33.09342, 31.42733,
  41.34376, 41.63763, 39.75784, 38.98249, 39.26605, 38.83189, 39.65921,
    38.46698, 35.43023, 35.16776, 35.46698, 36.18555, 36.48527, 36.17438,
    36.42402, 36.22709, 35.6164, 35.7401, 35.83401, 35.81164, 37.37441,
    37.91948, 36.89205, 35.53888, 35.10822, 35.189, 35.62875, 37.76955,
    36.03972, 32.24276,
  38.62775, 37.73642, 38.41263, 39.70662, 40.85919, 42.08347, 40.6528,
    36.75642, 34.85513, 35.07698, 34.62107, 34.51583, 34.66627, 35.29771,
    36.53222, 37.18892, 37.35836, 37.77358, 36.75073, 35.59332, 35.738,
    35.24171, 34.1922, 33.62676, 33.84196, 34.3443, 34.50113, 34.55306,
    35.12878, 32.83878,
  38.0643, 37.95957, 38.24712, 38.18777, 38.78793, 41.67698, 42.03743,
    37.37804, 35.01914, 35.7539, 36.41374, 36.93457, 37.2719, 37.98431,
    38.53485, 38.58438, 37.61319, 36.37097, 35.39825, 34.14194, 33.41985,
    33.2005, 33.02151, 32.90049, 33.00272, 33.60076, 33.64494, 33.06424,
    32.64037, 31.75678,
  22.1452, 22.18679, 22.21763, 22.24043, 22.23528, 22.22707, 22.23148,
    22.25263, 22.3238, 22.39399, 23.2039, 23.2434, 22.37857, 22.57035,
    22.66822, 22.34565, 22.24959, 22.28334, 22.31194, 22.807, 23.06255,
    22.62663, 22.58019, 23.04907, 23.27787, 22.92877, 25.29199, 26.90259,
    24.24732, 22.89537,
  22.45661, 22.48617, 22.34554, 22.59094, 22.43258, 22.28421, 22.33481,
    22.39615, 22.48517, 22.63624, 23.0052, 23.47201, 23.72202, 23.13483,
    22.87711, 22.86187, 22.40238, 22.44395, 22.8816, 23.33319, 23.27989,
    22.76415, 22.78669, 23.4517, 27.31024, 27.89697, 26.12094, 29.12415,
    25.03909, 23.47188,
  22.3888, 22.41249, 22.39115, 22.44898, 22.41056, 22.36969, 22.38497,
    22.45158, 22.53844, 22.59304, 22.69075, 23.04122, 23.29092, 23.67961,
    23.72246, 23.01017, 22.92748, 23.26089, 23.34107, 23.53766, 24.26173,
    25.43331, 26.3392, 25.91246, 30.4344, 32.82711, 28.40374, 28.62494,
    24.89419, 23.99474,
  22.41114, 22.4282, 22.57902, 22.72067, 22.97099, 23.40084, 23.42893,
    23.21345, 23.29094, 23.48267, 23.50224, 23.88596, 23.72237, 23.32137,
    24.15981, 24.96029, 24.31826, 23.49785, 23.69688, 24.075, 26.33117,
    27.58811, 26.75762, 31.19679, 32.91631, 30.03283, 30.74512, 27.89736,
    24.73403, 23.30941,
  22.85201, 22.68089, 22.92035, 23.24475, 23.47689, 23.65994, 23.71449,
    23.55364, 24.01764, 24.27323, 24.09924, 24.09895, 23.94911, 24.13065,
    24.70147, 25.16498, 24.41036, 23.8334, 24.28675, 28.51107, 29.838,
    25.72723, 25.64006, 27.8107, 29.74586, 29.11514, 27.85487, 28.436,
    28.94701, 24.71916,
  23.0176, 23.13909, 23.85443, 24.75486, 24.53446, 24.09946, 24.33587,
    24.15111, 23.78805, 23.80623, 23.81559, 25.53106, 27.51691, 27.62316,
    26.97311, 33.10647, 38.9617, 31.80098, 26.99125, 28.92215, 27.37907,
    24.45486, 25.04184, 26.00004, 28.78503, 28.27866, 30.60674, 41.73316,
    37.77069, 24.28162,
  23.5421, 23.86143, 24.61173, 25.44466, 25.36568, 25.09292, 26.07436,
    27.53008, 27.64254, 27.62736, 28.34054, 27.99409, 27.07669, 27.16776,
    31.67635, 38.1063, 36.06706, 29.20295, 26.74677, 26.54675, 25.24196,
    24.41465, 25.08258, 27.61787, 29.16463, 26.90623, 35.51812, 48.73466,
    37.51111, 22.96293,
  24.50892, 24.90299, 25.78354, 26.72617, 26.61505, 28.5715, 30.79577,
    28.86946, 27.38231, 27.45205, 27.44211, 26.51333, 25.56299, 25.68173,
    27.68558, 29.22089, 28.21385, 26.88535, 25.47877, 25.12148, 24.57263,
    24.39059, 25.83344, 28.37293, 27.98832, 26.47159, 38.38814, 42.94923,
    28.80816, 23.12152,
  27.31662, 27.67178, 28.69193, 28.9367, 29.67909, 31.35594, 30.12218,
    28.35954, 28.03495, 27.76101, 27.0302, 26.01954, 25.36451, 28.41052,
    30.21414, 27.27088, 27.09116, 28.56275, 28.54418, 26.27945, 24.51293,
    26.06108, 30.37598, 30.98079, 27.59203, 28.16356, 34.65408, 33.09391,
    25.08972, 23.10223,
  31.50086, 33.1018, 34.58965, 35.88022, 36.16679, 32.95889, 29.00041,
    28.28428, 27.40231, 26.41477, 27.24017, 30.62407, 32.00581, 31.17921,
    29.70107, 29.6821, 30.48061, 31.01838, 29.62088, 28.15748, 28.19608,
    29.16677, 30.31999, 28.84423, 33.53023, 41.93806, 35.79944, 26.10876,
    23.59318, 22.42496,
  43.6701, 46.7281, 43.75435, 39.14081, 37.93436, 35.85421, 32.15062,
    33.51567, 34.14692, 40.60201, 43.59843, 31.6457, 28.50132, 27.9155,
    27.2391, 28.08712, 29.32924, 29.4098, 28.32982, 28.19944, 30.57513,
    30.40452, 27.53905, 25.73451, 29.72388, 33.45886, 28.01195, 23.18404,
    22.76042, 22.2796,
  57.60332, 48.98376, 50.84565, 51.99973, 49.50171, 43.40486, 45.27333,
    41.7338, 35.17588, 39.07478, 38.49031, 26.77483, 27.7965, 28.62702,
    27.06094, 27.51682, 27.1739, 27.225, 26.74286, 27.24773, 30.10242,
    29.17246, 25.39042, 28.60731, 30.29613, 25.01119, 22.74638, 23.06685,
    22.98271, 22.45463,
  68.13518, 64.82087, 77.8422, 82.56182, 80.11588, 70.57519, 55.66282,
    39.45513, 35.68294, 33.5792, 30.65129, 25.41616, 30.14522, 32.16052,
    28.45857, 27.79943, 27.94921, 27.23416, 26.52356, 28.55294, 30.18371,
    27.63391, 25.11704, 29.89474, 30.97111, 24.32376, 22.91599, 23.26461,
    23.48436, 22.70024,
  75.57758, 101.1916, 99.48434, 95.57427, 85.95068, 73.75035, 60.95494,
    55.62296, 45.04874, 40.81581, 45.7186, 45.31004, 48.83581, 48.83,
    42.42212, 33.74355, 28.48196, 29.81447, 30.9891, 31.90944, 29.5914,
    28.84744, 30.29086, 27.56175, 25.26447, 23.58975, 22.99281, 22.83293,
    23.21307, 22.67896,
  58.25858, 66.35968, 64.13808, 61.42577, 54.89642, 57.15033, 73.60679,
    71.93595, 60.45737, 59.48938, 56.69473, 44.98167, 37.53529, 43.02811,
    43.88802, 32.26695, 31.48062, 31.83381, 34.58007, 35.3737, 32.12782,
    29.53798, 26.79597, 24.248, 23.29309, 23.67478, 23.08446, 22.68596,
    22.70544, 22.44079,
  46.0916, 45.7034, 44.72855, 42.92113, 41.58879, 45.77967, 52.69239,
    50.27227, 46.1708, 44.0903, 40.89183, 33.5649, 29.58412, 33.7173,
    33.58881, 31.11681, 32.48438, 31.31674, 32.37117, 31.9987, 27.76333,
    25.4971, 23.38932, 23.21434, 23.65208, 23.60325, 23.1589, 22.76391,
    22.62308, 22.36879,
  43.41335, 41.79066, 40.14763, 39.36665, 40.01189, 40.35322, 39.89444,
    38.74782, 36.65285, 34.29262, 30.44626, 30.27785, 33.6557, 32.30555,
    31.14607, 31.25443, 30.89377, 29.36033, 30.7733, 29.41906, 24.17879,
    24.31673, 23.90678, 23.40052, 23.40161, 23.58788, 23.08716, 22.55451,
    22.51108, 22.34601,
  39.50214, 38.58175, 37.75597, 38.23153, 38.46262, 38.57698, 37.75961,
    36.34751, 34.50238, 30.95282, 30.17045, 33.20679, 34.00225, 33.46901,
    34.73864, 32.86083, 29.0977, 27.1264, 29.81825, 28.49221, 24.31597,
    24.64269, 24.30844, 23.68687, 23.08852, 23.22466, 22.88428, 22.39061,
    22.36416, 22.28092,
  38.96457, 38.93565, 37.79089, 37.35183, 37.29183, 36.54966, 35.3401,
    33.68736, 31.2736, 29.28598, 31.61652, 32.37541, 29.29282, 29.97023,
    30.53143, 29.54495, 29.18534, 29.83743, 32.27615, 30.89894, 27.02169,
    25.31467, 24.36702, 23.83458, 23.01968, 22.88545, 22.72713, 22.39099,
    22.3292, 22.25694,
  39.65914, 39.62791, 37.99038, 36.53552, 36.26394, 35.33847, 33.94412,
    32.20787, 30.34942, 31.26971, 32.23464, 29.02014, 27.02503, 27.09283,
    26.62516, 25.99877, 27.44198, 29.75563, 31.61826, 32.02057, 30.03304,
    26.91144, 24.61454, 24.04582, 23.37685, 22.90191, 22.67973, 22.43428,
    22.34332, 22.26358,
  39.30708, 39.32259, 37.54417, 36.03248, 35.51982, 34.89423, 33.67788,
    32.04667, 31.05461, 32.00163, 29.98851, 26.16403, 26.33725, 26.49514,
    25.89255, 25.32109, 25.82862, 26.77526, 28.08278, 28.54977, 28.47089,
    27.91304, 26.31361, 24.72471, 23.71739, 23.10216, 22.65998, 22.42414,
    22.35671, 22.27297,
  39.6258, 38.66453, 37.11117, 36.14785, 35.70268, 34.88573, 33.91132,
    32.28463, 31.80128, 31.08288, 27.27268, 24.84046, 25.55133, 25.74133,
    25.55595, 25.42199, 25.16672, 25.17109, 25.54294, 25.50754, 26.51034,
    26.79953, 26.44796, 26.66941, 25.32179, 23.51749, 22.75614, 22.5277,
    22.37699, 22.27962,
  39.27885, 38.60479, 36.82929, 35.97843, 36.50562, 36.55075, 35.23152,
    32.73746, 31.60427, 29.22694, 25.36757, 24.47427, 25.0537, 25.29996,
    25.11004, 25.4763, 25.31313, 24.51595, 24.27473, 24.29193, 25.26892,
    25.1981, 24.66609, 26.29428, 26.69395, 24.38942, 22.93921, 22.92896,
    22.64224, 22.30461,
  38.73582, 38.30864, 37.59699, 37.49018, 37.70175, 37.37735, 36.54935,
    34.64903, 33.10338, 28.88736, 24.97898, 25.10568, 25.79418, 26.27128,
    26.13022, 26.24587, 26.25888, 25.29862, 24.38749, 24.35466, 24.50628,
    24.34075, 24.12169, 24.60477, 25.8656, 25.86251, 24.29984, 23.24666,
    22.94368, 22.4216,
  38.92388, 39.79794, 37.75798, 37.17581, 37.4657, 36.94513, 35.63445,
    34.20127, 33.75966, 29.44064, 25.23739, 25.60653, 26.31393, 26.67549,
    26.79881, 26.8592, 26.43939, 25.98813, 25.07184, 24.3285, 24.41087,
    24.46719, 24.3784, 23.9172, 23.91942, 25.19101, 25.21525, 23.97189,
    23.75927, 22.7684,
  39.49317, 41.73214, 40.20423, 38.41234, 37.18715, 35.9616, 35.92775,
    35.66087, 33.09464, 28.57698, 25.9215, 26.28127, 27.01101, 26.75085,
    26.28997, 26.33785, 26.01243, 25.83822, 25.37501, 24.62243, 24.84616,
    24.93669, 24.11953, 23.53681, 23.55448, 24.18765, 25.38824, 24.5928,
    23.7159, 22.67233,
  40.46017, 42.43055, 39.89841, 37.83782, 36.72789, 35.42245, 36.0629,
    35.46474, 31.08763, 27.17963, 26.25093, 26.58116, 26.82694, 26.46691,
    26.10168, 25.86484, 25.55359, 25.62212, 25.28143, 24.59278, 25.07821,
    26.11814, 26.01802, 25.16797, 24.98621, 25.08991, 26.69253, 26.33571,
    23.63024, 22.21922,
  39.95474, 40.67332, 38.52003, 37.53145, 37.74551, 36.98959, 36.69146,
    33.85895, 28.89309, 26.56112, 25.93093, 26.17197, 26.30741, 26.21017,
    26.4486, 26.18233, 25.49707, 25.41841, 25.70636, 25.9566, 26.80017,
    26.91992, 26.24937, 25.48916, 25.47056, 25.52542, 25.9138, 27.74219,
    26.1643, 22.88062,
  37.28767, 36.78264, 37.23541, 38.36739, 39.39407, 40.05433, 37.78529,
    32.34221, 28.13834, 26.35013, 25.02486, 24.69701, 24.87964, 25.32178,
    26.17699, 26.60676, 26.58584, 26.88846, 26.40078, 25.8021, 25.89651,
    25.42895, 24.5127, 24.07941, 24.34287, 24.80205, 24.85601, 24.9728,
    25.62743, 23.40498,
  35.97099, 36.07857, 36.41177, 36.61504, 37.23536, 39.36545, 38.37115,
    32.11117, 27.68082, 26.47861, 26.12516, 26.45542, 26.87439, 27.22551,
    27.52839, 27.71791, 26.91834, 25.99509, 25.45375, 24.54345, 23.97298,
    23.82049, 23.57447, 23.44856, 23.55107, 24.07127, 24.12697, 23.60328,
    23.30302, 22.50937,
  14.08992, 14.11846, 14.15515, 14.18215, 14.16153, 14.14125, 14.149,
    14.17348, 14.22188, 14.23935, 15.02139, 15.01868, 14.26211, 14.4987,
    14.58139, 14.27289, 14.20363, 14.23395, 14.24527, 14.7307, 14.9439,
    14.53898, 14.48975, 14.8878, 15.01694, 14.6756, 17.05293, 18.32978,
    15.93273, 14.70504,
  14.40714, 14.38556, 14.3034, 14.53834, 14.35143, 14.20037, 14.23428,
    14.28071, 14.34959, 14.47391, 14.89529, 15.36675, 15.58063, 15.02288,
    14.83673, 14.77435, 14.33363, 14.37333, 14.79304, 15.24108, 15.17004,
    14.59872, 14.5591, 15.16498, 18.77665, 18.86289, 18.23548, 21.01452,
    16.94863, 15.31615,
  14.35738, 14.34974, 14.33109, 14.40032, 14.30478, 14.22188, 14.23996,
    14.3007, 14.39849, 14.45976, 14.53251, 14.9075, 15.21482, 15.60367,
    15.59716, 14.85781, 14.77653, 15.04914, 15.05711, 15.18833, 15.75216,
    16.77383, 17.63076, 17.10596, 21.85077, 23.95387, 20.31844, 20.66285,
    16.83737, 15.82685,
  14.30791, 14.28582, 14.46261, 14.58397, 14.76291, 15.1354, 15.14613,
    14.95914, 15.04333, 15.23457, 15.25112, 15.62318, 15.397, 15.13625,
    15.93367, 16.65284, 15.97425, 15.07944, 15.06506, 15.226, 17.48083,
    18.72907, 18.13749, 22.14211, 23.46963, 21.77165, 22.83329, 20.00861,
    16.70967, 15.23348,
  14.68464, 14.43485, 14.65205, 14.98276, 15.24728, 15.40084, 15.36681,
    15.19704, 15.78125, 16.19517, 16.09509, 15.89639, 15.52596, 15.63617,
    16.21889, 16.60157, 15.67933, 14.98126, 15.2803, 19.44436, 20.71984,
    17.18161, 17.15696, 19.37247, 20.9122, 20.45728, 19.77279, 20.34745,
    20.50462, 16.35463,
  14.6363, 14.65975, 15.38293, 16.39734, 16.38166, 15.87235, 15.8535,
    15.64727, 15.3979, 15.4716, 15.36039, 16.90478, 18.53736, 18.51673,
    17.78168, 23.57667, 28.5352, 21.9391, 17.85773, 20.19345, 18.87997,
    15.99103, 16.55915, 17.32775, 19.97019, 19.36661, 21.44773, 31.62732,
    28.1578, 16.0004,
  14.70262, 15.00554, 15.85165, 16.81908, 16.93906, 16.50026, 17.14919,
    18.63529, 18.87665, 18.8176, 19.45064, 19.06734, 18.10896, 17.96862,
    22.52123, 29.16413, 27.24706, 20.32347, 18.07, 17.92604, 16.71474,
    15.94019, 16.47383, 18.73042, 20.22203, 17.78824, 26.36029, 39.61008,
    28.88642, 14.78244,
  14.88763, 15.20943, 16.1272, 17.03945, 16.95271, 18.93057, 21.01113,
    19.32144, 18.20731, 18.46028, 18.58136, 17.49107, 16.40562, 16.5025,
    19.1329, 21.03979, 19.6818, 18.07745, 16.85653, 16.58233, 16.13393,
    15.97302, 17.17456, 19.52863, 19.21939, 17.26972, 29.65445, 34.55,
    20.46367, 14.91104,
  16.22474, 16.40808, 17.44551, 17.63553, 18.28722, 20.44902, 19.81848,
    18.0846, 18.17801, 18.42015, 17.85906, 16.83403, 16.27613, 19.36493,
    20.95719, 18.23302, 18.20656, 19.5162, 19.41381, 17.47337, 15.95193,
    17.16319, 20.93162, 21.57735, 18.65295, 18.71907, 25.27038, 24.1573,
    16.59714, 14.93345,
  18.52538, 19.73907, 21.35539, 22.62165, 23.09861, 20.46083, 17.36178,
    17.16656, 17.10583, 16.5841, 17.77673, 20.97306, 22.21463, 21.91318,
    20.91418, 20.70329, 21.27845, 21.80492, 20.95646, 19.83885, 19.65845,
    20.67993, 21.88128, 20.3841, 24.49686, 32.23106, 26.68137, 17.804,
    15.48064, 14.3253,
  27.42311, 30.07136, 28.1981, 24.36994, 23.74854, 22.62126, 19.81218,
    21.46039, 23.10882, 29.53802, 32.10023, 22.6859, 19.99647, 19.4723,
    18.82883, 19.74212, 21.03627, 21.20188, 20.24322, 20.17375, 22.45135,
    22.41097, 19.59984, 17.67812, 21.71074, 25.75132, 20.39232, 15.20426,
    14.64207, 14.16999,
  39.56922, 31.78182, 33.51114, 34.56442, 32.63211, 28.64255, 31.25702,
    29.14635, 24.75063, 29.6972, 28.98181, 18.34643, 19.2114, 20.21052,
    18.97739, 19.40607, 19.15509, 19.2672, 18.85365, 19.34585, 22.18421,
    21.16268, 17.29973, 20.44239, 22.27201, 17.12776, 14.67569, 14.92036,
    14.87478, 14.3546,
  45.82278, 43.60081, 59.34008, 64.10822, 62.55853, 54.73046, 41.83122,
    28.27752, 25.99819, 24.78993, 21.30574, 16.39795, 21.33752, 23.77802,
    20.22129, 19.61075, 19.79912, 19.07071, 18.52776, 20.83311, 22.53167,
    19.62365, 16.92832, 22.08965, 23.37922, 16.32797, 14.79342, 15.13648,
    15.35985, 14.60726,
  56.56181, 79.32234, 81.15873, 76.20838, 66.82472, 57.50414, 48.44189,
    42.46578, 34.08821, 30.95738, 35.4806, 35.6784, 40.30523, 40.67166,
    33.87149, 25.2735, 20.09493, 21.486, 23.00971, 24.09328, 21.71218,
    21.01447, 22.68008, 19.96351, 17.44765, 15.46738, 14.8965, 14.74666,
    15.1222, 14.59984,
  44.58513, 53.32793, 51.8573, 49.10769, 42.85028, 45.53715, 60.14927,
    58.46238, 48.78013, 49.64584, 48.84621, 37.28522, 29.86108, 35.35401,
    36.04364, 23.98508, 22.93123, 23.17863, 25.23884, 26.53682, 24.552,
    22.10245, 19.61277, 16.6105, 15.05902, 15.47445, 14.98395, 14.59675,
    14.63226, 14.36463,
  33.706, 34.05884, 33.86686, 32.74911, 31.53368, 36.46953, 43.76952,
    40.97744, 37.7615, 37.36971, 33.8085, 25.75178, 21.19304, 25.67197,
    25.70642, 22.77865, 24.26937, 22.73134, 23.03942, 23.27563, 20.24666,
    17.94219, 15.66062, 15.44343, 15.61063, 15.39121, 15.00508, 14.70098,
    14.55509, 14.28527,
  31.842, 31.05282, 29.79308, 29.01929, 29.49146, 30.31819, 30.53967,
    29.42162, 27.99168, 26.21389, 22.12293, 22.12394, 24.90629, 23.41221,
    22.90813, 23.08295, 22.92408, 20.99558, 21.71877, 20.76921, 16.21012,
    16.30464, 16.05261, 15.6728, 15.47578, 15.42542, 14.93124, 14.48636,
    14.46468, 14.27481,
  29.03619, 28.24496, 27.20754, 27.57081, 28.06726, 28.74285, 28.7684,
    27.98578, 26.34101, 23.07626, 21.89639, 24.83807, 25.77868, 25.01575,
    26.62908, 25.00878, 21.2443, 18.99835, 21.18547, 19.98952, 16.22085,
    16.5007, 16.25402, 15.76989, 15.08783, 15.10705, 14.78461, 14.30597,
    14.28926, 14.20059,
  28.51652, 28.36968, 27.11406, 26.92163, 27.38421, 27.53894, 27.28296,
    26.17554, 23.7844, 21.51787, 23.2565, 24.1694, 21.56797, 22.30951,
    23.08086, 22.06005, 21.36014, 21.59956, 23.2218, 21.70362, 18.56974,
    17.13131, 16.23862, 15.77546, 14.92627, 14.76714, 14.63383, 14.30844,
    14.24705, 14.17548,
  29.00126, 29.07555, 27.63, 26.59821, 26.86321, 26.7049, 26.11675, 24.81897,
    22.83081, 23.28661, 24.14541, 21.22948, 19.27694, 19.30978, 18.91716,
    18.47868, 19.73388, 21.71159, 22.64815, 22.63365, 21.41296, 18.74185,
    16.40991, 15.92349, 15.27745, 14.8035, 14.59386, 14.33923, 14.24787,
    14.17703,
  28.74797, 29.11974, 27.66677, 26.49862, 26.39754, 26.29796, 25.70864,
    24.46948, 23.42889, 24.39654, 22.62953, 18.69558, 18.7369, 18.60091,
    17.85068, 17.36807, 17.84384, 18.68743, 19.47462, 19.78364, 20.24715,
    19.89981, 18.03458, 16.59816, 15.72503, 15.04378, 14.57169, 14.32699,
    14.24883, 14.17725,
  29.38079, 28.97466, 27.61615, 26.80511, 26.5505, 26.07015, 25.71203,
    24.67267, 24.41057, 24.07188, 20.33384, 17.29067, 17.75848, 17.72496,
    17.38126, 17.24633, 17.04529, 16.99698, 17.3892, 17.47128, 18.66682,
    18.78382, 17.96804, 18.302, 17.13223, 15.41705, 14.65703, 14.41531,
    14.27423, 14.18652,
  29.47095, 29.2092, 27.4721, 26.65403, 27.16649, 27.5048, 27.06518,
    25.34445, 24.58816, 22.53629, 18.41071, 16.79331, 17.10345, 17.24042,
    16.97653, 17.31611, 17.19407, 16.44304, 16.30435, 16.36265, 17.52014,
    17.24355, 16.26832, 17.87918, 18.31781, 16.23984, 14.89107, 14.84246,
    14.54253, 14.21304,
  29.14376, 28.95888, 28.09367, 28.03322, 28.45833, 28.62972, 28.74548,
    27.67651, 26.23059, 21.93796, 17.73358, 17.28793, 17.72211, 18.06868,
    17.85264, 17.97709, 18.032, 17.11942, 16.2999, 16.34483, 16.50412,
    16.2384, 15.90533, 16.29257, 17.36816, 17.59548, 16.24946, 15.18098,
    14.85806, 14.32286,
  29.40625, 30.23707, 28.39858, 27.99595, 28.59409, 28.54976, 27.97601,
    27.11934, 26.61399, 22.27325, 17.85101, 17.62881, 18.03302, 18.39948,
    18.45312, 18.38718, 18.01266, 17.65923, 16.91996, 16.34048, 16.23986,
    16.19818, 16.20835, 15.81935, 15.80239, 17.20716, 17.32197, 15.95097,
    15.69166, 14.71033,
  30.01159, 32.4536, 30.94429, 29.2112, 28.50119, 27.64586, 27.92774,
    28.02608, 25.80141, 21.55583, 18.51155, 18.20214, 18.58094, 18.43565,
    18.01838, 17.91877, 17.56955, 17.45437, 17.19641, 16.63692, 16.63139,
    16.6296, 15.99566, 15.54986, 15.57157, 16.25202, 17.5255, 16.63036,
    15.74412, 14.69045,
  31.40974, 34.02937, 31.38683, 29.01813, 27.94333, 26.82873, 28.13358,
    28.15345, 24.14207, 20.23743, 18.87272, 18.61193, 18.55538, 18.19548,
    17.76029, 17.47698, 17.17171, 17.18777, 17.07721, 16.60679, 16.8376,
    17.796, 17.76007, 17.11259, 17.03123, 17.13523, 18.81462, 18.34151,
    15.65658, 14.24099,
  31.56269, 32.81788, 29.9586, 28.3559, 28.50291, 27.88712, 28.29324,
    26.5341, 22.20186, 19.61794, 18.57026, 18.20382, 17.97587, 17.90013,
    18.02405, 17.71965, 17.05926, 16.9338, 17.47481, 18.00472, 18.52775,
    18.5462, 18.01306, 17.48255, 17.61526, 17.59853, 18.05255, 19.85722,
    18.14596, 14.81374,
  29.05394, 28.29735, 28.34641, 29.46538, 30.08269, 30.37954, 29.22339,
    25.15513, 21.43687, 19.35364, 17.52107, 16.76469, 16.81488, 17.0999,
    17.7017, 17.99809, 17.90113, 18.15979, 18.10317, 17.89248, 17.922,
    17.41246, 16.5025, 16.11124, 16.43186, 16.86969, 16.91191, 17.10275,
    17.73557, 15.39049,
  27.33203, 27.16556, 27.54399, 28.00841, 28.43611, 30.2653, 29.8706,
    24.81516, 20.75201, 19.16387, 18.18811, 18.23804, 18.72924, 18.82063,
    18.86995, 19.05612, 18.33732, 17.54094, 17.22421, 16.53219, 15.99834,
    15.85963, 15.57719, 15.42977, 15.53911, 16.09584, 16.26771, 15.67508,
    15.30527, 14.47108,
  13.68166, 13.70661, 13.73187, 13.7553, 13.75353, 13.74475, 13.7494,
    13.75622, 13.79928, 13.81463, 14.48566, 14.50937, 13.82629, 14.01465,
    14.10599, 13.85289, 13.79385, 13.80942, 13.79345, 14.22554, 14.44187,
    14.05266, 13.98574, 14.3589, 14.44782, 14.06377, 16.14605, 17.41465,
    15.3796, 14.29368,
  13.97069, 13.9647, 13.85625, 14.08132, 13.93573, 13.7965, 13.8189,
    13.85729, 13.91056, 14.02629, 14.46517, 14.89042, 15.01538, 14.51073,
    14.35631, 14.30862, 13.90726, 13.9195, 14.26877, 14.71293, 14.68782,
    14.11572, 14.00012, 14.49744, 17.58266, 17.71959, 17.49464, 20.33766,
    16.45398, 14.91447,
  13.95882, 13.95941, 13.91588, 13.9923, 13.89972, 13.79999, 13.80377,
    13.8734, 13.96122, 14.01571, 14.07555, 14.46167, 14.76734, 15.02067,
    14.99028, 14.35054, 14.24326, 14.48384, 14.50656, 14.59839, 15.01546,
    15.84281, 16.62714, 16.05738, 20.51654, 22.86234, 19.55523, 20.1019,
    16.32571, 15.42072,
  13.88823, 13.87203, 14.02374, 14.11334, 14.26858, 14.60223, 14.60521,
    14.42403, 14.47592, 14.6395, 14.66291, 15.03155, 14.83297, 14.5838,
    15.31881, 15.9778, 15.38116, 14.51911, 14.41917, 14.45296, 16.52444,
    17.76451, 17.12946, 20.77572, 22.29388, 21.02762, 22.1772, 19.41484,
    16.19507, 14.81477,
  14.18321, 13.97083, 14.16252, 14.45854, 14.71984, 14.88983, 14.83878,
    14.62902, 15.13567, 15.58171, 15.55549, 15.32032, 14.90398, 14.98223,
    15.63303, 16.04836, 14.99409, 14.22716, 14.45125, 18.29449, 19.73675,
    16.50635, 16.35475, 18.57606, 19.99847, 19.56214, 19.21366, 19.68813,
    19.67428, 15.77955,
  14.13356, 14.11248, 14.78165, 15.73045, 15.7756, 15.30857, 15.27319,
    15.05124, 14.81893, 14.89557, 14.74274, 16.15624, 17.59649, 17.55415,
    16.83941, 21.96467, 26.41236, 20.54124, 16.87134, 19.27428, 18.20028,
    15.38962, 15.92865, 16.56277, 18.95562, 18.44396, 20.27573, 30.51725,
    27.59885, 15.48735,
  14.14894, 14.41536, 15.23203, 16.18441, 16.36222, 15.83645, 16.23945,
    17.57192, 17.7176, 17.60499, 18.15515, 18.01679, 17.27974, 16.97745,
    21.08688, 27.6027, 26.18592, 19.54397, 17.38273, 17.29099, 16.11348,
    15.37463, 15.82951, 17.84209, 19.3148, 16.92912, 25.14071, 39.29571,
    29.15243, 14.31345,
  14.3094, 14.61824, 15.47388, 16.3061, 16.15591, 17.82697, 19.77294,
    18.35163, 17.27129, 17.49064, 17.68112, 16.63369, 15.54787, 15.5396,
    18.28687, 20.41674, 18.99769, 17.36366, 16.273, 16.06605, 15.6386,
    15.40277, 16.42922, 18.70399, 18.58641, 16.48917, 29.04855, 34.84529,
    20.35537, 14.48976,
  15.41036, 15.54336, 16.46385, 16.57591, 17.11022, 19.40711, 18.97248,
    17.13338, 17.18681, 17.43982, 16.9061, 15.87646, 15.31056, 18.41172,
    20.01365, 17.43737, 17.5335, 18.79041, 18.60728, 16.82344, 15.37437,
    16.44931, 20.08895, 20.83156, 18.01564, 17.91435, 24.79007, 23.97303,
    16.03942, 14.56043,
  17.3145, 18.27235, 19.77643, 21.16175, 21.68148, 19.26434, 16.33221,
    16.11743, 16.17038, 15.65708, 16.67376, 19.62351, 20.93094, 20.96779,
    20.13626, 19.74048, 20.20665, 20.7661, 20.12769, 19.10953, 18.96289,
    20.14244, 21.49671, 20.01556, 23.73271, 31.32706, 26.30333, 17.517,
    15.0868, 13.93214,
  24.13284, 26.54732, 25.36595, 22.10698, 21.85863, 20.85876, 18.19744,
    19.80804, 21.13846, 27.05674, 29.88388, 21.75057, 19.36595, 18.79726,
    18.08809, 18.99804, 20.19249, 20.32777, 19.4658, 19.49789, 21.88854,
    22.06283, 19.31272, 17.2899, 21.4052, 25.77192, 20.45685, 14.88818,
    14.22716, 13.76102,
  33.45201, 26.67925, 28.4792, 29.4009, 27.90095, 24.64371, 27.68606,
    26.44049, 22.7897, 27.81368, 27.61061, 17.81711, 18.46019, 19.3829,
    18.29743, 18.68364, 18.40403, 18.49223, 18.1487, 18.79282, 21.82512,
    20.84347, 16.92022, 19.93242, 21.90666, 16.93793, 14.33115, 14.47389,
    14.41797, 13.93198,
  42.18232, 37.00487, 46.50299, 52.82006, 52.12178, 46.62616, 36.32298,
    24.80573, 23.87663, 23.12041, 20.04472, 15.83159, 20.51824, 22.8209,
    19.45033, 18.82611, 19.03654, 18.28765, 17.83487, 20.28222, 22.17159,
    19.28713, 16.62257, 21.90173, 23.36711, 15.99635, 14.34267, 14.68876,
    14.88419, 14.18511,
  49.46407, 67.37472, 69.34579, 68.95502, 63.93957, 53.86647, 40.30067,
    36.65356, 29.58121, 26.96919, 32.04206, 33.11404, 38.03151, 38.72568,
    32.25818, 24.18704, 19.43766, 20.76863, 22.4221, 23.65041, 21.33837,
    20.4883, 22.18932, 19.85669, 17.31179, 15.04999, 14.44711, 14.31206,
    14.68848, 14.20474,
  35.67991, 43.76004, 44.38436, 44.32542, 39.39555, 39.3527, 50.16904,
    49.78535, 40.35954, 42.29449, 43.80667, 34.88858, 28.95022, 34.10326,
    34.4693, 23.19687, 22.38645, 22.6167, 24.37182, 25.76305, 23.85319,
    21.58081, 19.37027, 16.2958, 14.57314, 14.995, 14.51706, 14.17608,
    14.22779, 13.97191,
  24.83781, 25.41118, 26.17577, 25.67387, 23.83345, 28.14048, 35.67089,
    33.15693, 31.09808, 32.83269, 31.22788, 24.4838, 20.47003, 24.79331,
    24.75886, 22.12689, 23.79795, 22.20081, 22.2353, 22.62159, 19.76935,
    17.56005, 15.2631, 14.97086, 15.14155, 14.92548, 14.55043, 14.28153,
    14.14277, 13.88615,
  23.36798, 22.74523, 21.78795, 20.89352, 20.95425, 22.03102, 22.98815,
    22.7346, 23.06297, 23.20128, 20.46429, 20.98882, 23.78163, 22.43121,
    22.20031, 22.54458, 22.62061, 20.5379, 21.10477, 20.32092, 15.77336,
    15.79526, 15.49339, 15.17044, 15.02316, 14.97951, 14.50022, 14.07598,
    14.04422, 13.87074,
  20.92376, 20.08632, 19.04181, 19.19654, 19.68623, 20.54286, 21.30332,
    21.78773, 21.60057, 20.0166, 19.87944, 23.46198, 24.94221, 24.36217,
    26.23765, 24.80569, 21.15495, 18.54101, 20.63102, 19.49802, 15.58807,
    15.82481, 15.62556, 15.24599, 14.65553, 14.65836, 14.36868, 13.90723,
    13.88002, 13.79429,
  20.49422, 20.10977, 18.7547, 18.47587, 18.9675, 19.42305, 19.80155,
    19.76375, 18.9181, 18.32827, 21.23753, 23.06785, 21.1334, 22.1165,
    23.09043, 22.04601, 21.06576, 20.68299, 22.36299, 21.00684, 17.76722,
    16.44635, 15.64134, 15.24912, 14.48561, 14.33363, 14.21496, 13.89454,
    13.82699, 13.76247,
  20.92786, 20.71291, 19.21183, 18.16374, 18.42892, 18.43169, 18.35284,
    18.16065, 17.87695, 20.06711, 22.30251, 20.44811, 18.97051, 19.13717,
    18.78443, 18.27054, 19.31371, 20.86303, 21.75092, 21.98397, 20.69595,
    18.09133, 15.85853, 15.4289, 14.8263, 14.36683, 14.16868, 13.91633,
    13.82729, 13.76563,
  20.51456, 20.6126, 19.20263, 18.05008, 17.93629, 17.89168, 17.77418,
    17.7625, 18.49442, 21.29788, 21.09583, 18.1358, 18.49705, 18.35887,
    17.47498, 16.89202, 17.26169, 17.9791, 18.79072, 19.26018, 19.79779,
    19.30259, 17.34024, 16.13556, 15.32658, 14.63176, 14.1562, 13.91482,
    13.83688, 13.77284,
  20.95353, 20.34719, 19.05461, 18.23959, 17.96881, 17.61323, 17.7784,
    18.06506, 19.57145, 21.16913, 19.11004, 16.79166, 17.44109, 17.3588,
    16.89324, 16.67562, 16.49307, 16.48987, 16.94241, 16.99931, 18.12868,
    18.28865, 17.44761, 17.74207, 16.59229, 14.95083, 14.23312, 14.02732,
    13.86283, 13.76809,
  21.06392, 20.45143, 18.81834, 18.03244, 18.51993, 18.95743, 19.15295,
    18.79453, 19.84826, 19.87415, 17.29024, 16.21524, 16.64852, 16.71461,
    16.46385, 16.81238, 16.68747, 16.01232, 15.90646, 15.92029, 16.9879,
    16.74556, 15.8092, 17.3394, 17.69062, 15.69383, 14.45772, 14.42543,
    14.11137, 13.80342,
  20.76011, 20.25281, 19.33545, 19.26069, 19.81611, 20.26321, 21.08484,
    21.29605, 21.47532, 19.10873, 16.44843, 16.57269, 17.13794, 17.54466,
    17.35532, 17.45456, 17.44077, 16.55375, 15.86432, 15.97933, 16.10946,
    15.7518, 15.36903, 15.76952, 16.82801, 17.03017, 15.776, 14.77582,
    14.43976, 13.9156,
  20.81124, 20.97975, 19.59009, 19.48168, 20.38473, 20.81404, 20.73848,
    20.77941, 21.65519, 19.22544, 16.34167, 16.85717, 17.54621, 17.97176,
    17.98581, 17.87103, 17.47805, 17.09086, 16.42851, 15.96141, 15.80187,
    15.68346, 15.67304, 15.30778, 15.36323, 16.79688, 16.91959, 15.58802,
    15.29962, 14.31315,
  21.24479, 22.73144, 21.93652, 20.91356, 20.6463, 20.28863, 20.70523,
    21.39222, 20.63553, 18.51681, 16.89139, 17.36764, 18.06678, 17.97236,
    17.48856, 17.38218, 17.05385, 16.91009, 16.66722, 16.17521, 16.15094,
    16.08635, 15.44987, 15.02119, 15.07285, 15.83373, 17.17592, 16.30619,
    15.37155, 14.31746,
  22.61845, 24.34706, 22.68565, 21.08492, 20.09712, 19.22662, 20.98823,
    21.81089, 19.16774, 17.35806, 17.41009, 17.81649, 17.96973, 17.60654,
    17.1392, 16.89216, 16.64462, 16.67879, 16.57764, 16.13131, 16.28406,
    17.11772, 17.05161, 16.4345, 16.40282, 16.58923, 18.35019, 17.91969,
    15.21788, 13.83409,
  23.29648, 24.06436, 21.52939, 20.37539, 20.41062, 19.8988, 20.92739,
    20.16588, 17.42886, 16.87428, 17.22275, 17.46686, 17.36182, 17.23638,
    17.381, 17.12129, 16.53035, 16.43176, 16.97056, 17.53374, 17.85503,
    17.79661, 17.36036, 16.88561, 17.04674, 17.07284, 17.6404, 19.47318,
    17.74428, 14.40863,
  21.43234, 20.42632, 20.40822, 21.63708, 21.96462, 21.97445, 21.33422,
    18.54241, 16.74117, 16.73452, 16.31707, 16.11351, 16.23627, 16.53519,
    17.15299, 17.41548, 17.32788, 17.59951, 17.59484, 17.45145, 17.40336,
    16.86762, 16.00188, 15.62279, 15.97419, 16.43704, 16.56281, 16.89331,
    17.46525, 15.03498,
  20.27072, 19.84764, 20.2505, 20.82434, 21.07167, 22.39572, 22.07424,
    18.53166, 16.51091, 16.76883, 16.95582, 17.40393, 17.88528, 17.9995,
    18.17602, 18.39653, 17.70835, 17.00216, 16.75346, 16.10218, 15.56414,
    15.40678, 15.12922, 14.99309, 15.12738, 15.72285, 15.95387, 15.38604,
    14.98713, 14.09863,
  10.85241, 10.8737, 10.90869, 10.92383, 10.92622, 10.93034, 10.93035,
    10.93918, 10.97388, 10.98085, 11.67536, 11.75836, 11.01471, 11.1873,
    11.3055, 11.03439, 10.96592, 10.9894, 10.97434, 11.42118, 11.68867,
    11.30125, 11.22829, 11.60012, 11.63512, 11.20573, 13.34433, 14.85742,
    12.69839, 11.56662,
  11.17015, 11.18337, 11.05132, 11.28167, 11.12854, 10.98772, 11.01141,
    11.03026, 11.08723, 11.22707, 11.72987, 12.19941, 12.30029, 11.80109,
    11.60866, 11.56378, 11.10458, 11.11224, 11.48142, 12.02445, 12.05,
    11.37272, 11.19103, 11.6736, 14.85041, 15.43865, 14.91244, 18.32684,
    13.96382, 12.30477,
  11.18809, 11.19544, 11.13976, 11.23372, 11.10175, 10.98171, 10.97458,
    11.04007, 11.14624, 11.22395, 11.29978, 11.72798, 12.12373, 12.42484,
    12.36884, 11.61253, 11.46788, 11.76188, 11.79067, 11.89442, 12.27288,
    13.11011, 13.8702, 13.09334, 18.01384, 21.56525, 17.24838, 18.255,
    13.87277, 12.88391,
  11.10541, 11.08176, 11.25523, 11.34385, 11.46609, 11.80067, 11.80152,
    11.61852, 11.679, 11.86706, 11.9467, 12.32452, 12.13361, 11.93605,
    12.71318, 13.38052, 12.80083, 11.82921, 11.65754, 11.5727, 13.67924,
    15.15676, 14.35665, 18.42277, 20.79824, 19.05224, 20.41316, 17.48592,
    13.7552, 12.22451,
  11.45562, 11.18047, 11.37913, 11.67058, 12.00312, 12.17835, 12.0455,
    11.83521, 12.39967, 13.01947, 13.03435, 12.69257, 12.1705, 12.29449,
    13.05723, 13.52503, 12.34143, 11.31926, 11.47938, 15.52921, 17.40616,
    13.78541, 13.55784, 16.22319, 17.9507, 17.29626, 17.15657, 17.48984,
    17.33929, 13.1857,
  11.36488, 11.26373, 11.93286, 12.98118, 13.18657, 12.66473, 12.49695,
    12.27605, 12.10581, 12.3112, 12.13716, 13.36635, 14.87707, 14.94616,
    14.22088, 19.28793, 24.33351, 18.27249, 14.13054, 16.86298, 15.89872,
    12.58967, 13.1908, 13.91917, 16.45856, 16.17828, 17.51618, 28.36582,
    26.15149, 12.90733,
  11.28671, 11.54657, 12.43582, 13.54003, 13.88871, 13.29282, 13.52805,
    14.8735, 15.01097, 14.92734, 15.50141, 15.44978, 14.6845, 14.28415,
    18.57529, 25.95663, 24.74241, 17.28445, 14.88979, 14.88318, 13.53589,
    12.65914, 13.1339, 15.2506, 16.93423, 14.40306, 22.63027, 38.27734,
    28.14233, 11.60869,
  11.42309, 11.76196, 12.70736, 13.63716, 13.55274, 15.15192, 17.17142,
    15.78324, 14.63375, 14.8967, 15.12572, 14.03134, 12.71007, 12.62006,
    15.75966, 18.53186, 16.81622, 14.82868, 13.73501, 13.5657, 13.0364,
    12.71381, 13.79903, 16.21723, 16.16977, 13.87305, 26.99551, 34.37304,
    18.37057, 11.77788,
  12.56616, 12.69495, 13.70233, 13.8776, 14.34848, 16.91303, 16.59505,
    14.38789, 14.36549, 14.71012, 14.1066, 12.93139, 12.26406, 15.59966,
    17.74705, 15.01543, 15.03878, 16.56273, 16.44363, 14.45819, 12.67506,
    13.76341, 17.5737, 18.56379, 15.46118, 15.32995, 22.92442, 22.65162,
    13.44325, 11.86928,
  14.77618, 15.6128, 17.12197, 18.8491, 19.34948, 16.88359, 13.70429,
    13.32444, 13.25986, 12.65311, 13.57776, 16.78374, 18.2982, 18.58784,
    17.93654, 17.47248, 17.99386, 18.71681, 18.15701, 16.82714, 16.49087,
    17.77415, 19.32618, 17.78335, 21.40935, 29.94032, 25.23052, 15.31919,
    12.45077, 11.14395,
  20.69897, 23.78817, 23.19146, 19.79178, 19.46304, 18.58971, 15.90098,
    17.45679, 18.43901, 24.10158, 27.68834, 19.34955, 16.96196, 16.45945,
    15.7568, 16.76717, 18.13756, 18.33026, 17.38774, 17.23712, 19.79185,
    20.02025, 17.07655, 14.79692, 19.22825, 24.43833, 18.91765, 12.27558,
    11.46869, 10.9223,
  34.61942, 27.23747, 25.85532, 27.07389, 25.52327, 22.10407, 25.59119,
    24.68383, 20.48994, 25.61757, 25.96049, 15.27044, 16.02135, 17.20163,
    16.11411, 16.52238, 16.15787, 16.26269, 15.94121, 16.62603, 19.91513,
    18.86006, 14.4044, 17.532, 20.1008, 14.80935, 11.68047, 11.71588,
    11.64013, 11.11378,
  48.33704, 37.56681, 43.38676, 50.73891, 51.09678, 46.57452, 36.26142,
    23.06576, 22.08601, 21.5147, 18.45359, 13.03442, 18.21018, 21.24485,
    17.35279, 16.58701, 16.80856, 16.03942, 15.65088, 18.52987, 20.68689,
    17.13213, 14.08544, 19.96989, 22.02647, 13.51332, 11.5943, 11.9437,
    12.1473, 11.42316,
  52.03654, 67.16002, 68.01246, 69.60033, 64.50941, 54.36911, 40.75835,
    36.5336, 29.22022, 25.41057, 30.50411, 31.19433, 36.50285, 36.73923,
    30.65686, 22.72771, 17.42608, 19.05709, 20.8682, 22.39771, 19.76884,
    18.47794, 20.67401, 18.11544, 15.12996, 12.33356, 11.71547, 11.57377,
    11.97597, 11.4601,
  35.04996, 42.61774, 43.68801, 44.86111, 40.35111, 39.58107, 50.87845,
    50.98432, 39.75547, 40.68498, 42.3879, 33.75059, 27.0333, 32.15738,
    33.68452, 21.61873, 20.75, 21.13684, 23.06718, 24.70655, 22.49564,
    19.94816, 17.69298, 14.13289, 11.81169, 12.25997, 11.76095, 11.41373,
    11.47236, 11.19412,
  23.86568, 24.50167, 25.8569, 25.59371, 23.8537, 28.25481, 36.16148,
    33.06295, 30.29136, 31.88234, 30.28736, 23.2056, 18.60086, 23.32819,
    23.41797, 20.40734, 22.28672, 20.63057, 20.6051, 21.26574, 18.07524,
    15.50724, 12.86679, 12.53191, 12.52449, 12.16139, 11.78178, 11.52127,
    11.3658, 11.08599,
  22.68604, 22.28057, 21.53548, 20.53875, 20.49604, 21.86977, 23.04977,
    22.46098, 22.66702, 22.82279, 19.51405, 19.51633, 22.30079, 20.60631,
    20.63963, 21.17931, 21.19047, 18.7786, 19.18014, 18.68563, 13.44164,
    13.26536, 13.00773, 12.75592, 12.41684, 12.20149, 11.71947, 11.31205,
    11.27305, 11.07522,
  20.31468, 19.68919, 18.61605, 18.72994, 19.30847, 20.35395, 21.18325,
    21.55228, 21.09935, 19.11259, 18.40297, 22.05686, 23.51292, 22.65741,
    25.46037, 24.00866, 19.66799, 16.33138, 18.53689, 17.65292, 13.08393,
    13.32931, 13.09384, 12.73199, 12.00019, 11.93011, 11.64145, 11.11021,
    11.08987, 10.99164,
  20.03601, 19.70557, 18.2523, 17.95871, 18.52847, 19.11832, 19.55076,
    19.45379, 18.36713, 17.22168, 19.74637, 21.54381, 19.21849, 20.46261,
    22.19826, 20.92851, 19.37499, 18.33744, 20.26441, 19.11139, 15.51422,
    14.09008, 13.0737, 12.64246, 11.78679, 11.57907, 11.48516, 11.12205,
    11.02373, 10.94807,
  20.51691, 20.28658, 18.74566, 17.63064, 17.94053, 18.02375, 18.02448,
    17.80596, 17.22624, 19.09007, 21.14228, 18.77857, 16.94436, 17.29351,
    17.15604, 16.52197, 17.45078, 18.94077, 19.86607, 20.1093, 18.62543,
    15.89865, 13.30401, 12.8021, 12.16001, 11.6244, 11.41371, 11.14012,
    11.02054, 10.95113,
  20.09323, 20.20475, 18.75536, 17.54644, 17.48487, 17.53004, 17.4438,
    17.36474, 17.93813, 20.59334, 20.09919, 16.41524, 16.57501, 16.35813,
    15.39294, 14.7504, 15.15745, 15.91098, 16.6667, 17.14933, 17.74634,
    17.21397, 14.88048, 13.58756, 12.70782, 11.94421, 11.41346, 11.13882,
    11.03401, 10.95651,
  20.69136, 19.97902, 18.66323, 17.85631, 17.62941, 17.28706, 17.50598,
    17.77193, 19.26908, 20.74285, 18.13789, 15.09331, 15.48812, 15.21655,
    14.61051, 14.33165, 14.10718, 14.10262, 14.59073, 14.65981, 16.0064,
    16.25356, 15.06737, 15.3871, 14.11691, 12.32327, 11.46926, 11.22845,
    11.04982, 10.95613,
  20.9535, 20.25498, 18.52013, 17.70303, 18.24138, 18.79474, 19.11312,
    18.74964, 19.78816, 19.57671, 16.24275, 14.48604, 14.55739, 14.41578,
    14.00038, 14.32654, 14.28022, 13.61559, 13.47655, 13.46714, 14.76653,
    14.5972, 13.3001, 15.0249, 15.40852, 13.17292, 11.72187, 11.69571,
    11.33198, 10.98113,
  20.7268, 20.15141, 19.09279, 19.00081, 19.68997, 20.33846, 21.45215,
    21.93101, 21.98856, 18.87466, 15.20192, 14.70151, 14.82043, 15.02573,
    14.79312, 14.97623, 15.10884, 14.17394, 13.34339, 13.49586, 13.80906,
    13.37073, 12.79931, 13.29295, 14.49444, 14.64159, 13.20027, 12.13935,
    11.73404, 11.12149,
  20.63382, 20.67407, 19.33763, 19.38369, 20.58165, 21.35663, 21.49118,
    21.69299, 22.34979, 18.99478, 14.94659, 14.81169, 15.09531, 15.42308,
    15.49047, 15.5244, 15.20377, 14.71918, 13.93839, 13.48143, 13.37092,
    13.19692, 13.15607, 12.76184, 12.78438, 14.298, 14.50529, 13.0532,
    12.6685, 11.60893,
  20.95057, 22.186, 21.74619, 21.21761, 21.16677, 21.11285, 21.76259,
    22.38186, 20.98033, 18.00156, 15.29438, 15.22302, 15.70252, 15.56141,
    15.07019, 15.03415, 14.72123, 14.55, 14.30024, 13.72086, 13.68479,
    13.64847, 12.94489, 12.39866, 12.37544, 13.20526, 14.68305, 13.79793,
    12.7696, 11.65958,
  22.26867, 23.66096, 22.75799, 21.72435, 20.81602, 20.00108, 22.00769,
    22.61277, 19.12636, 16.47551, 15.75619, 15.74185, 15.73172, 15.23959,
    14.70854, 14.46023, 14.2216, 14.29068, 14.20361, 13.64153, 13.80224,
    14.77741, 14.71236, 13.93986, 13.82104, 14.05798, 15.97158, 15.55271,
    12.61971, 11.10064,
  23.46343, 24.12004, 21.65354, 21.00359, 21.01999, 20.47404, 21.50226,
    20.50299, 17.06563, 15.88375, 15.64241, 15.43367, 15.07848, 14.83147,
    14.96984, 14.66348, 14.02359, 13.983, 14.50836, 15.0513, 15.51865,
    15.63972, 15.13062, 14.46727, 14.56738, 14.64497, 15.32935, 17.26442,
    15.46243, 11.74748,
  22.00212, 20.99393, 20.76759, 22.22208, 22.58907, 22.6067, 21.87414,
    18.71159, 16.37405, 15.86468, 14.73475, 13.94943, 13.75171, 13.97876,
    14.6892, 14.94459, 14.81967, 15.17424, 15.1709, 15.03133, 15.07751,
    14.54239, 13.55476, 13.05653, 13.43947, 13.96731, 14.11324, 14.53072,
    15.20373, 12.50463,
  20.83402, 20.40192, 20.74355, 21.22974, 21.56251, 22.99023, 22.59761,
    18.67468, 16.07763, 15.798, 15.23558, 15.09061, 15.3101, 15.51332,
    15.8253, 16.00952, 15.30913, 14.54087, 14.17198, 13.49646, 12.97412,
    12.79934, 12.48998, 12.33721, 12.49359, 13.1182, 13.41012, 12.82377,
    12.37407, 11.37864,
  12.22318, 12.24418, 12.27767, 12.29449, 12.29695, 12.29346, 12.30729,
    12.34184, 12.37165, 12.37746, 13.12106, 13.24456, 12.40124, 12.56477,
    12.71949, 12.42729, 12.33798, 12.36162, 12.3501, 12.82402, 13.15191,
    12.73842, 12.65366, 13.04048, 13.05045, 12.58712, 14.82286, 16.56442,
    14.28174, 13.09325,
  12.51869, 12.5429, 12.39815, 12.64643, 12.51446, 12.36664, 12.40579,
    12.44703, 12.50496, 12.64771, 13.24037, 13.74578, 13.79014, 13.28405,
    13.0482, 13.00969, 12.49154, 12.49208, 12.90104, 13.53088, 13.59762,
    12.85261, 12.59977, 13.15753, 16.38157, 17.14704, 16.79697, 20.82375,
    15.87299, 13.9562,
  12.5755, 12.57928, 12.50985, 12.62687, 12.49472, 12.36933, 12.37653,
    12.44775, 12.56898, 12.66561, 12.739, 13.23453, 13.71824, 14.03529,
    13.98396, 13.0939, 12.85952, 13.22112, 13.2941, 13.41029, 13.72653,
    14.60815, 15.45691, 14.6846, 19.73409, 23.87504, 19.50588, 20.88562,
    15.80527, 14.62298,
  12.49973, 12.46736, 12.65481, 12.75171, 12.87716, 13.27846, 13.31046,
    13.07154, 13.09888, 13.28932, 13.39392, 13.83685, 13.68373, 13.49933,
    14.38049, 14.99996, 14.42059, 13.36839, 13.09182, 12.89575, 15.10494,
    16.94674, 16.10481, 20.3108, 23.06185, 21.5046, 23.48637, 20.05413,
    15.67765, 13.90215,
  12.91714, 12.58959, 12.80729, 13.09472, 13.43029, 13.70213, 13.62071,
    13.31817, 13.8553, 14.58294, 14.66926, 14.28661, 13.65319, 13.81286,
    14.79875, 15.28308, 13.86334, 12.61639, 12.72098, 16.8898, 19.35323,
    15.52507, 15.18768, 18.20621, 20.19925, 19.58123, 19.7245, 19.85257,
    19.54189, 14.92467,
  12.83103, 12.67031, 13.3722, 14.48943, 14.7046, 14.16434, 13.98024,
    13.73752, 13.60312, 13.86181, 13.6521, 14.90225, 16.71903, 16.99257,
    16.13563, 21.23845, 26.89321, 20.24349, 15.67779, 18.83748, 17.99726,
    14.10695, 14.78335, 15.69127, 18.52114, 18.35791, 19.36417, 31.38696,
    29.7016, 14.69786,
  12.67649, 12.93596, 13.93604, 15.19896, 15.5476, 14.86075, 14.98873,
    16.46988, 16.59707, 16.40962, 17.13393, 17.35398, 16.78627, 16.33868,
    20.91799, 29.5947, 28.39576, 19.49337, 16.77077, 16.87624, 15.2591,
    14.18079, 14.7474, 17.13199, 19.09175, 16.27572, 24.57591, 42.57786,
    32.63386, 13.20083,
  12.80848, 13.19826, 14.32076, 15.40222, 15.23109, 16.83932, 19.16801,
    17.82602, 16.42842, 16.68327, 17.12646, 16.01672, 14.39542, 14.15595,
    17.91493, 21.56575, 19.13724, 16.57051, 15.45909, 15.26991, 14.67119,
    14.28145, 15.46486, 18.20317, 18.2101, 15.50722, 30.11781, 39.85456,
    21.40987, 13.31111,
  14.02188, 14.25457, 15.40581, 15.57717, 15.97998, 19.15556, 19.08097,
    16.32041, 16.21342, 16.66891, 16.04962, 14.58141, 13.62714, 17.18622,
    19.90336, 16.94359, 16.76079, 18.48219, 18.36735, 16.27762, 14.2404,
    15.4182, 19.51362, 20.73162, 17.23458, 17.01957, 26.23184, 26.59862,
    15.27205, 13.45508,
  16.54209, 17.35979, 19.1732, 21.35796, 21.95282, 19.32866, 15.54922,
    15.04942, 15.1314, 14.44734, 15.16512, 18.55261, 20.30076, 20.93566,
    20.33724, 19.63272, 20.15809, 20.97118, 20.31715, 18.78397, 18.33374,
    19.71889, 21.59987, 19.95559, 23.68123, 33.32801, 28.57167, 17.53283,
    14.20842, 12.63213,
  22.16414, 25.89693, 25.50776, 21.9655, 21.74658, 21.12527, 18.12575,
    19.52794, 20.38266, 25.61913, 30.05124, 21.8904, 19.25647, 18.77709,
    17.87374, 18.971, 20.59402, 20.73269, 19.46114, 19.17244, 22.06011,
    22.46421, 19.25595, 16.63459, 21.81061, 28.32121, 22.08858, 13.995,
    12.97499, 12.31087,
  36.19219, 28.37791, 26.78345, 27.15845, 26.25162, 22.77723, 27.149,
    27.15056, 22.63372, 27.7475, 28.99841, 17.20951, 17.71806, 19.23014,
    18.26996, 18.77395, 18.30004, 18.34175, 17.82494, 18.57048, 22.41036,
    21.40046, 16.23705, 19.20262, 22.38913, 17.12727, 13.39043, 13.21569,
    13.10378, 12.52519,
  48.48986, 36.30897, 42.03368, 49.27026, 50.51582, 47.94925, 39.3203,
    24.43927, 24.01573, 24.35435, 20.69245, 14.4371, 19.9135, 23.5155,
    19.60154, 18.64183, 18.75719, 17.91791, 17.48236, 20.79282, 23.43718,
    19.30268, 15.78303, 22.04735, 24.90524, 15.58467, 13.06461, 13.43768,
    13.64247, 12.87927,
  53.21689, 60.43174, 62.20439, 64.9465, 62.72283, 56.83284, 44.41184,
    39.58131, 31.12293, 26.82096, 31.56266, 32.4678, 38.34473, 38.67324,
    33.62578, 24.91658, 19.37836, 21.07545, 23.23287, 25.22563, 22.40615,
    20.50684, 23.35252, 20.97709, 17.55766, 13.97597, 13.17796, 13.06727,
    13.49999, 12.93878,
  35.87315, 40.79557, 44.39848, 49.29602, 51.31326, 48.55301, 49.98035,
    51.67169, 39.61436, 40.18732, 43.64333, 36.18884, 29.66207, 34.65234,
    36.71618, 24.12633, 23.15379, 23.62265, 25.91783, 27.86135, 25.41245,
    22.91689, 20.81662, 16.55166, 13.35915, 13.82216, 13.25501, 12.88487,
    12.95894, 12.65394,
  23.81961, 26.31957, 30.07471, 32.08448, 31.42229, 31.96824, 35.54688,
    32.35648, 29.23076, 31.44651, 32.27079, 25.52484, 20.49524, 25.92147,
    26.11143, 22.84275, 25.11399, 23.40257, 23.28751, 24.38974, 21.09578,
    18.25079, 14.95206, 14.21769, 14.06721, 13.72113, 13.32397, 13.03327,
    12.85445, 12.52824,
  21.87194, 22.44434, 22.27678, 20.94389, 19.72995, 20.70063, 22.37545,
    21.55468, 21.96263, 23.05337, 20.58746, 20.82203, 24.11726, 22.62341,
    23.02726, 23.88646, 24.2702, 21.52763, 21.81791, 21.81607, 15.65336,
    15.1446, 14.72239, 14.48771, 14.07049, 13.78745, 13.26014, 12.81262,
    12.7477, 12.50947,
  18.74596, 18.13987, 16.83604, 16.53145, 16.96798, 18.25061, 19.22928,
    19.90467, 20.16338, 18.73161, 18.35682, 23.07465, 25.49776, 24.60098,
    28.43908, 27.44423, 22.7061, 18.82066, 21.2765, 20.57993, 14.95666,
    15.07708, 14.79932, 14.49295, 13.64449, 13.50876, 13.17969, 12.56267,
    12.52231, 12.40482,
  18.12387, 17.53736, 15.83429, 15.5034, 16.09491, 16.68917, 17.24112,
    17.45648, 16.76022, 15.98034, 19.46144, 22.5666, 20.81786, 22.68733,
    25.4534, 24.15683, 22.13174, 20.80462, 23.15641, 21.77028, 17.28108,
    15.88346, 14.85492, 14.38976, 13.36688, 13.11805, 13.00858, 12.55226,
    12.4409, 12.35539,
  18.46378, 17.86506, 16.19552, 14.97732, 15.29989, 15.44144, 15.55586,
    15.48227, 15.10952, 17.67522, 21.08261, 19.64653, 18.33103, 19.45313,
    19.82205, 19.18393, 20.14675, 21.74462, 22.76382, 22.87049, 20.82922,
    17.91585, 15.1188, 14.53187, 13.74928, 13.144, 12.90281, 12.58783,
    12.44325, 12.36042,
  17.85229, 17.653, 16.15331, 14.87755, 14.86117, 14.95849, 14.82136,
    14.69426, 15.65303, 19.51673, 20.35298, 17.22952, 18.26404, 18.68474,
    17.87731, 17.15976, 17.48757, 18.2415, 19.01829, 19.74637, 20.41049,
    19.62857, 16.82334, 15.36042, 14.30726, 13.49145, 12.91589, 12.58646,
    12.44683, 12.36463,
  18.45026, 17.38818, 16.05238, 15.24201, 15.04736, 14.578, 14.65687,
    14.9741, 17.21595, 20.00518, 18.34917, 15.99901, 17.41144, 17.59535,
    16.94164, 16.45717, 16.06695, 16.00424, 16.68008, 16.89502, 18.46477,
    18.83963, 17.10355, 17.41732, 15.92878, 13.91935, 12.95693, 12.67714,
    12.4711, 12.36307,
  18.73593, 17.71426, 15.94594, 15.06354, 15.58829, 15.99965, 16.28106,
    16.16223, 18.08119, 19.03125, 16.38925, 15.52413, 16.41462, 16.53,
    16.00847, 16.20534, 16.1472, 15.54035, 15.43651, 15.36316, 16.99108,
    16.95135, 15.12284, 17.14489, 17.45805, 14.85053, 13.18211, 13.15996,
    12.77783, 12.39464,
  18.5411, 17.71548, 16.50945, 16.25352, 16.96923, 17.70818, 19.10114,
    20.07293, 20.7985, 18.2916, 15.24181, 15.71356, 16.49008, 16.97133,
    16.69993, 16.89723, 17.11345, 16.08944, 15.075, 15.24037, 15.8438,
    15.35935, 14.5071, 15.19524, 16.50129, 16.46932, 14.81439, 13.6837,
    13.2446, 12.55956,
  18.47633, 18.25281, 16.6447, 16.58569, 18.03059, 19.2084, 19.74038,
    20.34164, 21.46654, 18.50677, 14.93767, 15.7517, 16.6737, 17.39676,
    17.57987, 17.69979, 17.29682, 16.62493, 15.68581, 15.21009, 15.16296,
    14.94208, 14.96037, 14.54892, 14.52288, 16.20388, 16.38131, 14.71886,
    14.27121, 13.11319,
  18.77862, 19.66082, 19.01609, 18.68814, 19.1091, 19.47882, 20.39901,
    21.31195, 20.08927, 17.3757, 15.17513, 16.02608, 17.22701, 17.54681,
    17.22542, 17.18846, 16.69548, 16.45756, 16.13721, 15.40897, 15.39629,
    15.40875, 14.67672, 14.02308, 13.94952, 14.93562, 16.57829, 15.59601,
    14.43276, 13.20036,
  20.12587, 21.19114, 20.41764, 19.63728, 19.08467, 18.50546, 20.96316,
    21.87697, 18.03734, 15.52914, 15.63827, 16.66399, 17.44463, 17.29468,
    16.79191, 16.47284, 16.15093, 16.2017, 16.04434, 15.30944, 15.45875,
    16.46119, 16.39202, 15.57024, 15.46803, 15.86032, 18.1196, 17.61854,
    14.27245, 12.56904,
  21.79469, 22.41686, 19.50917, 19.0647, 19.33002, 18.94923, 20.30541,
    19.3374, 15.48532, 14.795, 15.67312, 16.59088, 16.88777, 16.83849,
    17.01821, 16.68119, 15.91558, 15.75598, 16.21295, 16.68592, 17.21631,
    17.45774, 16.98393, 16.27533, 16.38503, 16.65749, 17.61764, 19.58737,
    17.42099, 13.26361,
  20.52815, 19.28529, 18.9561, 20.93772, 21.31212, 21.1672, 20.42418,
    16.9202, 14.49524, 14.83851, 14.86513, 15.05376, 15.3817, 15.85446,
    16.67659, 16.88435, 16.61364, 16.93946, 16.98297, 16.82497, 16.93062,
    16.40349, 15.29781, 14.75753, 15.21207, 15.84752, 16.05384, 16.59141,
    17.16654, 14.07888,
  19.62136, 19.00343, 19.56, 20.36873, 20.49832, 21.79553, 21.2301, 16.89936,
    14.43703, 15.1051, 15.5237, 16.17511, 16.8653, 17.29843, 17.70802,
    17.88086, 17.17347, 16.43987, 16.04433, 15.25613, 14.67543, 14.46904,
    14.09475, 13.9157, 14.13724, 14.83612, 15.0951, 14.40405, 13.96695,
    12.87077,
  17.9273, 17.9741, 18.00398, 18.02138, 18.02016, 18.01949, 18.02916,
    18.07614, 18.11277, 18.1497, 19.01462, 19.23171, 18.15545, 18.33529,
    18.55412, 18.20664, 18.0997, 18.12477, 18.1122, 18.64597, 19.0698,
    18.59942, 18.51147, 18.924, 18.94362, 18.47718, 20.93189, 23.37083,
    20.56299, 19.1517,
  18.21995, 18.28959, 18.11086, 18.40985, 18.24379, 18.08504, 18.13335,
    18.18968, 18.2673, 18.46584, 19.10051, 19.69846, 19.81198, 19.21356,
    18.8715, 18.91439, 18.2806, 18.28648, 18.80167, 19.511, 19.51951,
    18.67177, 18.36814, 19.1137, 22.77305, 24.57175, 23.6302, 29.07233,
    22.59945, 20.24526,
  18.2881, 18.31116, 18.24546, 18.36341, 18.22434, 18.09026, 18.10325,
    18.2091, 18.33789, 18.45, 18.57814, 19.11609, 19.64324, 20.03713,
    20.05051, 18.998, 18.74181, 19.2404, 19.27272, 19.3568, 19.81294,
    21.07247, 22.18215, 21.54987, 26.79185, 32.52776, 27.48483, 29.24751,
    22.53192, 21.08315,
  18.23416, 18.2035, 18.40753, 18.54505, 18.70989, 19.23894, 19.32826,
    19.01525, 19.00293, 19.17332, 19.3307, 19.85504, 19.71886, 19.38897,
    20.45707, 21.2612, 20.68546, 19.38822, 18.95541, 18.82456, 21.67927,
    24.24296, 23.11131, 28.02511, 31.40218, 29.08719, 32.68816, 28.12198,
    22.35167, 20.14637,
  18.7376, 18.30716, 18.56535, 18.94233, 19.37795, 19.72994, 19.67433,
    19.31552, 19.89079, 20.87952, 21.06606, 20.38882, 19.51896, 19.86153,
    20.94901, 21.32692, 19.88642, 18.42626, 18.72324, 24.00162, 27.52772,
    22.23912, 21.88286, 25.09233, 27.38499, 26.82276, 27.30866, 28.40373,
    28.06081, 21.57061,
  18.59643, 18.42796, 19.29972, 20.70023, 21.08311, 20.4416, 20.08914,
    19.82285, 19.58006, 19.83945, 19.62507, 21.04469, 23.36789, 23.58591,
    22.95498, 27.94545, 34.99302, 28.24166, 22.62267, 26.29891, 25.28086,
    20.32618, 21.12012, 22.31368, 25.34638, 25.48168, 26.11305, 40.59756,
    40.49327, 21.28095,
  18.46143, 18.82115, 20.04518, 21.56241, 22.13297, 21.36541, 21.17412,
    23.05776, 23.37416, 23.23237, 24.10884, 24.31124, 23.34326, 22.88873,
    27.70439, 36.61815, 35.59419, 26.68313, 23.51461, 23.61968, 21.68198,
    20.36584, 21.07515, 23.91906, 26.15491, 23.38233, 31.3492, 51.35321,
    42.83628, 19.58337,
  18.63023, 19.16021, 20.54412, 21.8796, 21.67878, 23.56278, 26.35946,
    24.6493, 22.91391, 23.34302, 23.85508, 22.56354, 20.51448, 20.44669,
    24.43406, 28.27677, 25.70156, 23.47187, 21.85137, 21.54434, 20.86135,
    20.40424, 21.93878, 25.20643, 25.21186, 22.77975, 37.66201, 49.55183,
    29.02666, 19.49984,
  20.29644, 20.63184, 21.787, 21.98883, 22.59179, 26.78931, 26.68487,
    22.74937, 22.79348, 23.32064, 22.57994, 20.78599, 19.75231, 23.92621,
    27.60629, 24.03862, 23.39993, 25.47139, 25.38164, 22.86691, 20.32062,
    21.88018, 26.75042, 28.32233, 24.05233, 24.41509, 34.3119, 35.4125,
    21.93902, 19.47404,
  22.98516, 23.62768, 26.12114, 29.6429, 29.93275, 26.82695, 21.94903,
    21.17471, 21.21758, 20.53638, 21.33115, 25.60818, 27.71203, 28.31526,
    27.38991, 26.49998, 27.23186, 28.26615, 27.46361, 25.47781, 25.0445,
    26.56353, 28.68619, 27.14703, 31.36821, 42.88581, 38.37932, 24.56393,
    20.2943, 18.45666,
  30.69206, 36.96254, 37.21075, 29.78057, 29.47665, 28.69227, 25.87607,
    26.98225, 28.26454, 33.31625, 39.40747, 29.60495, 26.46899, 25.80425,
    24.93766, 26.15091, 28.07554, 28.2869, 26.79378, 25.82108, 29.02047,
    29.51673, 25.98084, 23.10889, 28.8801, 36.11426, 29.39782, 19.92036,
    18.88799, 18.06424,
  47.19059, 38.60865, 35.6624, 33.3938, 33.43986, 28.22492, 33.4967,
    34.11721, 30.10367, 35.66576, 36.75818, 23.18881, 24.12943, 26.27946,
    25.16668, 26.01129, 25.46098, 25.44735, 24.67806, 25.37074, 29.8217,
    28.64863, 22.61106, 26.02522, 30.43202, 24.19107, 19.42365, 19.12705,
    19.01964, 18.33438,
  60.19814, 46.27232, 49.93996, 56.66348, 57.68716, 55.372, 49.63379,
    43.7649, 50.5012, 35.98604, 26.62697, 22.46629, 28.66748, 30.3022,
    27.35933, 25.7998, 26.03548, 24.89793, 23.99778, 27.61269, 30.95399,
    26.13446, 22.28448, 29.27116, 33.21857, 21.79086, 18.89274, 19.39699,
    19.63391, 18.77855,
  67.04805, 59.02151, 62.43295, 67.9334, 70.12125, 69.76936, 63.56649,
    62.87843, 51.39054, 35.76363, 39.70156, 42.37838, 48.23661, 48.80914,
    42.82759, 32.3014, 26.863, 28.81277, 31.3295, 33.6632, 30.29688,
    27.35691, 31.49806, 28.55307, 24.30232, 19.96596, 19.06845, 18.96374,
    19.41286, 18.83485,
  52.05716, 65.49017, 73.65117, 78.39595, 77.07889, 69.24906, 68.13445,
    69.07728, 47.96183, 48.83112, 56.93642, 49.17432, 42.23042, 44.54895,
    46.24163, 33.08513, 31.83231, 32.52698, 35.15819, 36.877, 32.68914,
    30.56602, 28.51877, 23.36873, 19.39973, 19.85616, 19.18544, 18.76811,
    18.77417, 18.46242,
  38.72879, 49.80747, 55.03433, 52.65743, 45.33881, 47.65863, 54.4735,
    40.39354, 43.8785, 52.44142, 41.27872, 35.69886, 30.84575, 35.20766,
    34.91525, 31.9585, 34.52027, 32.18389, 31.30514, 32.46927, 28.24652,
    25.19857, 21.59599, 20.416, 20.17314, 19.72608, 19.2448, 18.90106,
    18.62704, 18.28441,
  30.00189, 31.07037, 30.47425, 26.96083, 24.89771, 29.63997, 33.19537,
    28.57528, 34.30989, 36.74955, 26.21365, 27.0107, 31.77777, 30.28975,
    31.42389, 32.35007, 33.22036, 29.74146, 29.40772, 30.39357, 22.62826,
    21.60224, 20.86998, 20.57566, 20.0588, 19.7184, 19.18875, 18.64805,
    18.50451, 18.27891,
  23.45273, 22.81462, 20.77676, 20.16401, 21.20949, 23.11417, 24.17535,
    25.38175, 25.28503, 22.83596, 22.59742, 28.69942, 32.5769, 31.62181,
    37.55736, 36.46686, 31.1122, 26.17236, 29.06038, 28.69684, 21.2702,
    21.46793, 21.03012, 20.61608, 19.5423, 19.43111, 19.11338, 18.37062,
    18.29287, 18.1678,
  22.13474, 21.28517, 18.90218, 18.42144, 19.20809, 19.96032, 20.78363,
    20.88204, 19.70818, 18.56133, 22.94301, 27.64886, 26.30329, 29.2656,
    33.97466, 32.54636, 30.32055, 28.35674, 31.49078, 29.84595, 23.96305,
    22.43747, 21.21159, 20.59132, 19.31815, 19.02185, 18.90487, 18.3611,
    18.22506, 18.11617,
  21.91171, 20.90066, 18.84468, 17.33167, 17.79708, 18.0494, 18.18395,
    17.97068, 17.35844, 20.25264, 24.72456, 23.63119, 22.91505, 25.44909,
    26.89256, 26.68694, 28.03978, 30.11203, 31.0715, 31.07021, 28.10711,
    24.80694, 21.58844, 20.76267, 19.75703, 19.07434, 18.78649, 18.42075,
    18.21955, 18.11966,
  20.72528, 20.30317, 18.52775, 16.97968, 16.98555, 17.12675, 16.97498,
    16.69191, 17.70462, 22.24372, 23.72036, 20.4553, 22.7478, 24.38469,
    24.22972, 23.94323, 24.77535, 26.07598, 26.68754, 27.37131, 28.1173,
    27.3489, 23.49405, 21.70979, 20.29072, 19.47075, 18.80209, 18.42561,
    18.24407, 18.13737,
  21.48801, 19.77239, 18.24431, 17.27231, 17.11887, 16.50029, 16.5465,
    16.82418, 19.46651, 22.91306, 21.25289, 18.94269, 21.79171, 23.11965,
    23.15144, 23.05263, 22.92193, 22.98685, 23.80793, 24.05119, 25.65496,
    26.4002, 23.95309, 24.38093, 22.54745, 20.13178, 18.90185, 18.55089,
    18.25472, 18.13203,
  21.72285, 20.01653, 18.04016, 16.98052, 17.70426, 18.09076, 18.28835,
    18.1129, 20.42232, 21.82077, 18.77714, 18.41682, 20.63715, 21.87902,
    22.10147, 22.79407, 22.94067, 22.33225, 22.22616, 22.06867, 23.63855,
    23.97351, 21.88304, 24.35902, 24.63539, 21.38535, 19.17971, 19.11296,
    18.6173, 18.16963,
  21.42918, 19.87073, 18.74694, 18.39044, 19.19761, 19.82674, 21.64715,
    23.26685, 24.16374, 21.04921, 17.49727, 18.78147, 20.76533, 22.4338,
    22.93409, 23.54187, 24.04939, 23.02917, 21.78007, 21.93165, 22.68965,
    22.03924, 20.97037, 22.03125, 23.45344, 23.19237, 21.15882, 19.71569,
    19.1275, 18.37531,
  21.21894, 20.98732, 18.94334, 18.55746, 20.31879, 22.02582, 22.89743,
    23.85502, 24.93042, 21.51851, 17.2731, 18.98606, 21.0152, 22.96488,
    23.99057, 24.64879, 24.41429, 23.59255, 22.40325, 21.77728, 21.74564,
    21.36673, 21.49655, 21.16076, 20.90198, 22.67177, 22.78549, 20.81953,
    20.21874, 19.05691,
  21.8571, 23.01315, 21.85319, 21.22161, 21.83517, 22.69839, 24.17431,
    25.37313, 23.42019, 20.32448, 17.67445, 19.29301, 21.58305, 23.13327,
    23.6866, 24.23994, 23.74804, 23.26567, 22.79286, 21.78625, 21.77017,
    21.97437, 21.20933, 20.24293, 19.99501, 21.1687, 22.92798, 21.89498,
    20.44131, 19.18674,
  23.27221, 24.49934, 23.53762, 22.22522, 21.97609, 21.77458, 25.17077,
    26.41179, 21.20905, 18.06841, 18.18912, 19.92291, 21.7882, 22.83028,
    23.21164, 23.30177, 22.93985, 22.87101, 22.60686, 21.60536, 21.93787,
    23.24252, 23.08506, 21.83691, 21.62194, 22.17712, 24.63165, 24.37555,
    20.44569, 18.39666,
  25.84257, 27.48414, 22.153, 21.49492, 22.26793, 22.21875, 24.25125,
    23.31079, 18.16968, 17.07816, 18.20045, 19.87163, 21.23114, 22.35359,
    23.47274, 23.42806, 22.51241, 22.30745, 22.70378, 23.03844, 23.9376,
    24.5486, 23.8836, 22.79742, 22.69475, 23.17116, 24.30167, 26.58044,
    24.22433, 19.28514,
  24.16057, 22.49988, 21.63923, 25.54827, 25.62576, 24.52117, 24.21274,
    20.10143, 16.84369, 17.12263, 17.29845, 18.07197, 19.47328, 21.20155,
    23.03924, 23.63778, 23.30283, 23.66833, 23.6617, 23.3476, 23.66367,
    23.17102, 21.82503, 21.06072, 21.51928, 22.30324, 22.65359, 23.35028,
    23.80289, 20.33376,
  22.95431, 21.82892, 23.54997, 26.06728, 25.62196, 25.92824, 25.13695,
    20.01821, 16.81509, 17.55542, 18.05841, 19.33848, 21.20942, 22.8364,
    24.20243, 24.79061, 24.03407, 23.1596, 22.58598, 21.61249, 20.96557,
    20.67249, 20.24813, 20.02418, 20.32572, 21.14122, 21.4776, 20.73342,
    20.12039, 18.81888,
  28.45755, 28.57423, 28.65369, 28.69969, 28.67262, 28.6725, 28.70409,
    28.7691, 28.85481, 29.15829, 30.60857, 31.04502, 29.07256, 29.4567,
    29.83801, 29.09813, 28.86786, 28.92216, 28.96146, 29.796, 30.53628,
    30.14052, 30.5873, 31.55712, 32.34733, 32.79787, 36.76788, 40.39347,
    33.63125, 30.48283,
  29.1426, 29.39721, 28.99269, 29.53466, 29.16017, 28.82431, 28.9553,
    29.10551, 29.30246, 29.70923, 30.57347, 31.62339, 32.19338, 31.12186,
    30.26333, 30.45701, 29.33502, 29.58332, 30.58257, 31.60925, 31.52118,
    30.72041, 31.10852, 34.19376, 40.93789, 44.69522, 41.55556, 47.94228,
    35.85092, 31.99777,
  29.15939, 29.28644, 29.18997, 29.22875, 28.99352, 28.88153, 28.93649,
    29.14216, 29.37474, 29.53655, 29.8222, 30.72037, 31.57659, 32.40598,
    32.57763, 30.71246, 30.51028, 31.43916, 31.46558, 32.0641, 34.23023,
    38.18162, 40.66879, 41.34474, 49.40985, 56.13345, 48.51271, 47.83438,
    36.02487, 33.43502,
  29.14195, 29.22763, 29.58664, 29.92723, 30.31203, 31.23181, 31.35216,
    30.78163, 30.77573, 31.22569, 31.67564, 32.4143, 32.24119, 31.53827,
    33.59575, 35.26752, 34.19516, 31.78834, 32.01752, 33.95459, 40.46972,
    45.20359, 42.84, 50.1543, 56.50194, 51.12954, 55.98369, 46.00581,
    36.07383, 31.80754,
  30.15962, 29.48833, 30.08903, 30.79781, 31.52038, 31.89408, 31.76593,
    31.5087, 32.65431, 33.75501, 33.10938, 32.48034, 32.02485, 32.82901,
    34.40591, 35.0229, 33.52436, 31.99539, 34.90289, 43.46691, 48.46786,
    40.28996, 40.34895, 43.9872, 45.68086, 45.39763, 45.05609, 48.97152,
    45.93729, 33.28522,
  29.80493, 30.20504, 31.88421, 34.16928, 34.00163, 32.41513, 32.55682,
    31.87772, 31.33241, 31.53019, 31.91986, 35.62627, 40.7907, 40.15015,
    43.02177, 52.68056, 57.27615, 50.64865, 42.93065, 46.45365, 42.96589,
    35.91499, 37.71342, 40.50514, 43.80089, 46.64712, 52.7199, 66.86353,
    63.07647, 34.11617,
  29.76645, 31.06814, 33.18255, 35.31927, 34.953, 33.93208, 36.16429,
    39.63365, 40.15804, 40.11927, 41.99829, 41.82381, 39.82654, 41.53994,
    48.81365, 58.16157, 55.87524, 47.41028, 40.9121, 40.55394, 37.26032,
    35.30336, 37.44084, 43.05341, 47.82618, 49.27079, 58.55539, 72.15948,
    61.2482, 31.07535,
  29.3496, 30.95144, 33.44144, 35.45584, 35.08514, 39.16358, 45.85824,
    42.18664, 37.5034, 38.01923, 38.0262, 36.052, 34.29216, 36.27805,
    40.75395, 44.88516, 43.49058, 41.24157, 36.68368, 36.17678, 34.9766,
    35.11324, 39.14434, 45.16671, 46.88677, 48.37426, 62.74401, 70.10859,
    47.77658, 30.59721,
  31.02758, 31.64328, 34.41802, 35.66074, 36.68084, 41.98941, 40.47655,
    35.86514, 36.08686, 35.97992, 34.19468, 32.0973, 32.87133, 41.91376,
    48.92878, 41.55397, 40.02016, 43.25707, 43.32731, 39.13504, 35.84565,
    39.86553, 47.6067, 50.32119, 44.60132, 49.20702, 60.65899, 56.72892,
    36.95308, 30.5473,
  33.93109, 39.16624, 45.25185, 45.87634, 46.5255, 42.11847, 30.55972,
    30.20483, 29.4, 29.58757, 33.66652, 44.39014, 48.82763, 47.89534,
    44.53757, 45.2135, 47.4186, 47.68618, 45.17826, 41.3231, 42.64366,
    44.37149, 46.57679, 48.37387, 58.28909, 70.5865, 60.98129, 38.01575,
    31.37163, 29.01846,
  48.68695, 52.55854, 52.69906, 46.49729, 46.52697, 42.49981, 35.85609,
    39.58718, 45.14039, 52.99985, 57.79914, 43.77112, 39.50244, 39.43661,
    39.78544, 42.89736, 45.61319, 44.93388, 42.97026, 41.46995, 45.34783,
    45.9214, 41.29171, 39.50632, 46.16829, 51.00208, 41.17369, 30.09122,
    29.70347, 28.61486,
  64.88692, 50.08232, 50.99132, 53.64873, 53.2145, 45.04108, 52.54633,
    53.44012, 49.30994, 50.27341, 45.63713, 33.00426, 35.88496, 39.56386,
    40.55262, 42.68371, 42.07017, 41.61111, 40.65444, 42.31487, 46.01117,
    43.55429, 36.02192, 40.46203, 45.87076, 36.54512, 30.0258, 30.03283,
    29.8964, 28.98769,
  77.61427, 68.24712, 85.47507, 93.92405, 92.60502, 84.05913, 69.25834,
    52.20702, 52.93315, 42.33605, 35.55957, 32.373, 41.52513, 48.25418,
    46.43848, 42.58329, 43.22165, 41.49231, 40.62955, 48.05497, 50.08061,
    39.61287, 36.55857, 42.86007, 45.7728, 32.94524, 29.65314, 30.43331,
    30.64935, 29.59901,
  90.85725, 106.8363, 110.3991, 107.4548, 95.43081, 86.03039, 78.65836,
    72.3643, 57.72651, 50.50035, 61.63279, 64.03854, 70.14498, 72.17297,
    64.99435, 52.5363, 45.08656, 48.15235, 51.71428, 53.75578, 47.04913,
    40.67773, 46.43707, 40.47005, 34.47047, 31.07306, 30.00084, 29.78335,
    30.29246, 29.62582,
  89.83556, 89.30927, 86.44668, 78.77354, 68.74166, 70.16969, 85.3771,
    81.77897, 70.47982, 77.25713, 79.2157, 67.78674, 62.1124, 68.41963,
    67.52245, 54.96345, 54.93034, 57.47522, 61.41012, 60.33128, 50.39718,
    47.38878, 42.28802, 33.65561, 30.61284, 31.09079, 30.17916, 29.56965,
    29.49353, 29.0978,
  80.47799, 75.3189, 69.2142, 62.54866, 61.1059, 67.25348, 76.83371, 78.8792,
    78.21128, 64.69698, 63.74575, 53.99136, 49.06152, 56.83534, 56.85851,
    55.73933, 60.00003, 56.73512, 56.46361, 54.89969, 42.8917, 38.03617,
    33.63953, 31.46402, 31.43479, 30.92494, 30.20041, 29.67376, 29.29228,
    28.89001,
  62.1544, 55.93969, 50.2859, 49.02591, 50.62415, 52.53424, 58.93298,
    64.80655, 55.74083, 50.70693, 46.60084, 45.97992, 53.27045, 53.4548,
    54.95354, 56.68511, 56.3843, 50.44023, 50.56303, 49.55059, 34.5374,
    32.68642, 32.27232, 32.1146, 31.16601, 30.86285, 30.10098, 29.3068,
    29.14298, 28.883,
  44.71412, 41.16161, 38.62115, 40.4981, 43.70783, 47.84131, 50.37381,
    48.34958, 43.38483, 40.88676, 42.74409, 52.40301, 56.97, 58.92081,
    63.76421, 59.46709, 50.82712, 45.35577, 49.66068, 45.39171, 32.87444,
    34.29404, 33.49673, 32.27645, 30.35898, 30.36415, 29.99857, 28.96856,
    28.88146, 28.74275,
  39.96636, 38.89942, 35.88758, 35.89503, 40.43601, 42.8018, 40.64996,
    37.54374, 35.05993, 35.26934, 43.72414, 51.38322, 49.36212, 54.18573,
    55.67072, 49.80856, 49.01086, 52.58572, 55.53545, 49.21557, 38.93829,
    36.92258, 34.14596, 32.23601, 30.10445, 29.85215, 29.65459, 28.95991,
    28.78272, 28.66828,
  39.16253, 39.07662, 34.96621, 33.20083, 36.06213, 35.59977, 32.70451,
    30.99456, 31.09212, 39.1929, 48.37113, 45.10048, 43.81206, 45.73096,
    44.03704, 41.68077, 45.46445, 52.6976, 55.29191, 53.80085, 47.15893,
    40.16748, 34.63515, 32.49817, 30.75059, 29.9534, 29.52689, 29.06956,
    28.79083, 28.68012,
  37.92468, 37.52304, 33.102, 31.11403, 31.68648, 30.5847, 29.05745,
    29.36946, 33.64588, 43.48763, 45.84936, 38.64876, 40.62814, 40.10334,
    38.58445, 38.96714, 43.01497, 47.62844, 50.25508, 49.96096, 45.98414,
    41.98718, 37.45372, 33.73333, 31.42727, 30.53051, 29.56305, 29.08785,
    28.83503, 28.7072,
  38.71786, 36.06812, 31.76075, 30.17611, 29.61352, 27.95732, 28.69821,
    31.04012, 37.91063, 44.01262, 39.34248, 34.22006, 36.74986, 36.08945,
    36.14129, 38.68916, 42.12294, 44.52943, 45.38336, 43.60847, 41.66727,
    40.62818, 38.75003, 38.18468, 35.05505, 31.55846, 29.7455, 29.28702,
    28.86135, 28.72577,
  37.48297, 35.28653, 30.59052, 28.51856, 29.94803, 31.32113, 32.46881,
    33.57732, 38.92828, 40.78238, 32.85372, 30.55042, 32.10288, 33.20772,
    35.07315, 39.36341, 42.42323, 42.09522, 40.71484, 38.84531, 38.69955,
    38.48281, 36.91496, 39.08234, 38.73351, 33.66444, 30.13846, 30.0804,
    29.37114, 28.77971,
  37.16083, 34.59519, 32.64743, 31.85458, 33.30634, 34.98689, 37.64973,
    38.42878, 41.62056, 38.28568, 29.13547, 29.42538, 31.48333, 34.7489,
    38.07982, 41.66123, 43.77074, 41.814, 38.73874, 37.51811, 37.01856,
    36.37318, 36.02791, 37.07687, 38.0235, 36.62011, 33.14223, 30.83212,
    30.02745, 29.07501,
  35.78929, 37.20176, 32.0601, 31.58171, 34.70984, 36.44788, 37.59403,
    38.57201, 42.52452, 37.57815, 27.73009, 29.87024, 33.00417, 37.2362,
    40.80431, 43.5134, 43.47339, 41.56126, 38.19082, 35.63485, 35.90334,
    36.37012, 35.89721, 34.54724, 33.84247, 35.41384, 35.04839, 32.38062,
    31.48287, 30.0659,
  37.6791, 40.50273, 36.80931, 35.64974, 36.70109, 36.62568, 37.94438,
    40.40175, 41.00176, 34.35286, 29.02028, 32.10101, 35.92552, 38.79024,
    40.34815, 41.96479, 41.54473, 39.94497, 37.19271, 34.81391, 36.51913,
    37.3552, 34.49631, 31.96891, 31.7212, 33.21159, 35.20737, 34.03172,
    31.7222, 30.15565,
  41.10712, 44.05807, 40.79372, 38.06573, 37.74451, 36.08622, 38.57415,
    40.52789, 37.17376, 30.91077, 31.54682, 34.94743, 37.37554, 38.17823,
    38.73123, 39.65717, 39.4537, 38.2482, 36.1544, 34.4455, 36.59299,
    38.72321, 37.04288, 34.3272, 33.75119, 34.76999, 37.78463, 37.37063,
    31.79328, 29.04023,
  45.14808, 46.73839, 39.45784, 37.87196, 39.86819, 38.84282, 40.38752,
    38.77148, 32.2291, 30.84793, 33.62777, 36.20497, 36.85478, 36.91591,
    38.38623, 39.32235, 38.18059, 36.9518, 36.13943, 36.58194, 39.7335,
    40.93784, 38.14567, 35.7628, 35.20153, 36.23048, 37.70382, 40.25677,
    37.09269, 30.40955,
  40.27067, 35.57063, 36.12917, 40.72737, 42.82318, 44.79926, 42.57145,
    35.12469, 30.48412, 32.29731, 33.00484, 32.92599, 32.81919, 34.08354,
    37.22287, 39.39761, 39.61092, 39.55795, 38.02268, 37.1304, 38.55139,
    37.52712, 34.70055, 33.20963, 33.73993, 35.03584, 35.64919, 36.28397,
    36.29445, 31.88589,
  36.87989, 35.59919, 39.07621, 40.4393, 39.99432, 43.56533, 44.89829,
    36.07164, 31.54763, 33.65224, 34.1717, 34.55401, 35.31068, 36.99089,
    39.67822, 41.77942, 40.91619, 38.44027, 36.25286, 34.43117, 33.60033,
    32.7065, 31.94263, 31.62069, 32.14376, 33.25287, 33.64146, 32.72527,
    31.47469, 29.57843,
  36.23909, 36.65694, 37.11712, 37.58576, 37.80452, 38.17302, 38.68544,
    39.31183, 40.11884, 41.49406, 43.97341, 44.16841, 40.10922, 41.36997,
    42.14832, 41.30399, 42.17476, 44.20232, 46.65472, 50.23017, 52.58835,
    51.91803, 53.5926, 56.55597, 58.72047, 59.91077, 66.07927, 67.97961,
    47.46527, 41.16336,
  36.64725, 37.30898, 36.59352, 37.92755, 37.31744, 37.04542, 37.80925,
    38.51102, 39.48016, 40.79898, 42.81927, 45.42696, 47.04019, 44.97854,
    43.95754, 46.00631, 46.02673, 49.27872, 53.26614, 56.75869, 58.05651,
    58.74805, 61.10276, 67.20301, 73.27056, 70.37228, 64.93528, 69.17141,
    48.53001, 42.87092,
  33.31285, 33.59682, 34.10663, 34.59346, 34.94715, 35.4772, 36.04559,
    36.88541, 38.01612, 39.43504, 41.39225, 44.59688, 48.19717, 52.24006,
    54.93861, 54.05643, 57.43388, 62.0613, 65.63437, 71.14078, 78.77039,
    85.88132, 88.30598, 87.4034, 87.31878, 84.06441, 77.17332, 66.94573,
    49.39991, 45.00602,
  35.67652, 36.64867, 38.62254, 40.65786, 42.38729, 44.49942, 44.86438,
    44.44298, 45.70185, 47.68159, 49.72566, 52.53993, 55.068, 57.0832,
    64.23739, 69.17398, 68.11593, 66.87273, 72.71527, 79.53748, 89.74805,
    92.85481, 87.14081, 93.77528, 93.9741, 90.49293, 85.46893, 66.87731,
    50.70056, 42.74252,
  40.03319, 39.27173, 41.80606, 43.48518, 44.72945, 44.79826, 45.29287,
    46.42965, 49.53145, 52.30907, 52.93883, 55.94284, 59.07397, 62.94293,
    67.341, 70.71397, 70.51645, 68.44144, 73.88451, 83.61262, 86.77797,
    76.72453, 78.90828, 86.19202, 92.73673, 92.74273, 85.23951, 89.21654,
    78.33573, 50.98506,
  41.03991, 44.00404, 48.36564, 52.87083, 52.85922, 52.38327, 55.89586,
    58.54965, 60.54729, 65.48997, 72.72389, 85.07719, 96.63016, 94.69797,
    96.14599, 100.7496, 105.6884, 96.14448, 84.72524, 85.33479, 78.37029,
    72.1185, 78.06873, 84.47212, 91.21603, 89.88322, 84.62643, 97.70921,
    88.13441, 48.53527,
  47.9846, 54.1771, 61.03881, 68.31304, 72.73549, 78.75592, 88.61282,
    97.39293, 97.42957, 94.54963, 92.62476, 85.59616, 75.88211, 76.58996,
    78.99052, 82.90089, 83.96371, 79.7786, 72.65134, 74.2503, 72.00948,
    72.17884, 77.71776, 85.31837, 85.70506, 75.84026, 76.89755, 87.06258,
    74.68613, 40.99083,
  57.37354, 65.21043, 72.85965, 80.3187, 83.77359, 91.75613, 95.75662,
    77.96127, 66.14644, 64.80626, 60.26311, 55.57161, 52.70544, 55.60354,
    59.98185, 66.34875, 71.17193, 71.09924, 65.69437, 67.37894, 68.10667,
    71.44456, 78.95406, 83.8946, 78.66273, 73.82357, 82.49564, 82.46167,
    60.9978, 41.70116,
  68.89522, 72.80669, 76.87927, 78.12598, 76.67224, 78.38215, 68.33124,
    62.89864, 65.62318, 65.77268, 64.77827, 65.12885, 70.25975, 84.92682,
    94.12277, 79.93817, 81.8974, 88.40475, 88.19798, 81.56593, 79.57515,
    91.4719, 102.8924, 99.62279, 84.74277, 89.88435, 89.80046, 74.5337,
    48.34756, 41.11806,
  92.19897, 100.2663, 96.49583, 99.28522, 91.86801, 79.55914, 62.10917,
    70.93561, 74.55138, 83.89156, 95.08023, 107.792, 106.0068, 102.9077,
    98.49982, 105.8665, 109.7648, 107.9889, 101.4793, 98.78558, 105.3698,
    103.0252, 97.32076, 85.67271, 91.15932, 101.0719, 83.23103, 54.56212,
    40.8217, 37.99832,
  109.1494, 107.4483, 108.1241, 99.87514, 109.8634, 110.5735, 105.3674,
    110.367, 114.8356, 116.3048, 107.6661, 82.90315, 81.1937, 83.08305,
    86.87654, 92.47099, 96.36001, 95.37136, 92.11299, 91.60822, 100.9596,
    95.79969, 74.84193, 66.33244, 71.49823, 70.57201, 53.84297, 40.83783,
    39.91897, 37.81834,
  111.102, 105.1905, 111.4437, 113.1157, 114.488, 100.9478, 103.0007,
    97.05593, 87.96487, 76.90643, 71.22717, 68.92203, 76.2205, 82.26358,
    83.72826, 82.93571, 80.54698, 79.20334, 76.85561, 78.96857, 87.56574,
    80.73621, 63.36147, 71.10919, 73.53062, 55.4186, 40.72718, 42.41053,
    40.83562, 38.91477,
  118.9535, 119.1559, 122.0404, 122.9521, 121.6046, 117.2077, 106.8107,
    94.77103, 98.38847, 78.86212, 77.74966, 79.08691, 90.03371, 97.27132,
    91.52284, 78.28246, 79.10254, 76.21358, 74.90054, 80.97529, 83.8961,
    73.72949, 66.28384, 65.69954, 62.20985, 49.73774, 42.36515, 43.57133,
    42.67198, 40.27946,
  118.7255, 118.7396, 117.7197, 115.6809, 113.3222, 111.5482, 111.1182,
    111.4911, 109.309, 109.8227, 111.5243, 110.202, 113.2357, 114.8647,
    112.0439, 95.71207, 93.55997, 97.66791, 102.2231, 96.80209, 82.00716,
    70.34891, 66.41818, 54.32079, 47.95932, 45.62097, 42.60109, 41.39985,
    41.36115, 40.0109,
  104.7614, 98.0598, 101.8465, 105.9064, 108.5345, 110.2761, 114.398,
    115.3604, 113.089, 113.8871, 113.4594, 112.7638, 114.2174, 114.4457,
    113.328, 112.848, 109.4417, 106.4927, 104.9679, 93.16316, 68.82859,
    62.78878, 52.74686, 47.7279, 45.90694, 44.59515, 42.15686, 40.50943,
    39.49953, 38.72324,
  97.30721, 102.263, 107.9313, 110.5813, 111.3277, 113.5597, 116.0441,
    114.361, 112.9915, 113.275, 113.535, 111.6491, 107.868, 113.0731,
    112.4945, 107.7975, 103.7775, 91.09418, 84.54836, 73.40013, 54.70808,
    53.56108, 47.52571, 46.21705, 45.56459, 43.77789, 41.67672, 40.41713,
    39.26783, 38.49548,
  89.61442, 88.70866, 91.63045, 95.74409, 99.71877, 104.676, 109.1394,
    112.4091, 112.1612, 110.4969, 102.4928, 111.4717, 115.3142, 111.6234,
    104.6554, 95.71793, 86.92572, 77.79755, 76.01215, 70.06422, 51.40702,
    52.48266, 48.3345, 46.00502, 44.45382, 43.58644, 41.24816, 39.22449,
    38.79226, 38.41993,
  73.02545, 76.12527, 76.62961, 81.114, 85.55908, 91.49084, 96.09689,
    100.7115, 104.3594, 104.9915, 113.6707, 117.1955, 116.9952, 115.7913,
    112.5414, 93.47643, 75.27278, 70.33182, 76.90652, 70.11867, 53.20268,
    53.376, 49.12656, 46.87376, 43.35301, 42.1329, 40.7283, 38.43751,
    38.26892, 38.04211,
  78.66879, 76.10575, 69.04675, 67.91156, 73.64587, 78.95392, 85.15085,
    91.25579, 94.8764, 101.3598, 111.9524, 108.9776, 92.14516, 92.7287,
    89.3606, 84.36665, 87.53419, 94.03326, 96.13229, 82.70634, 61.76074,
    54.72219, 49.52232, 46.0864, 42.22638, 40.71785, 39.87505, 38.52689,
    38.12399, 37.9818,
  74.31012, 69.19911, 62.77125, 59.90407, 66.22809, 72.01108, 78.30803,
    83.58124, 89.32346, 98.54778, 98.77495, 79.58675, 75.62785, 76.40024,
    75.79774, 77.23679, 84.30821, 92.39238, 92.26607, 85.60292, 71.31754,
    58.78522, 50.38797, 46.67711, 43.69519, 41.16378, 39.94237, 38.76344,
    38.1363, 38.0309,
  65.5679, 61.92516, 57.2359, 56.82208, 62.43075, 67.75745, 72.0065,
    75.79639, 80.74676, 85.68679, 78.24605, 66.03864, 73.76506, 75.3165,
    74.3781, 73.31932, 75.21741, 76.26889, 76.01869, 72.39055, 67.07037,
    63.42562, 56.32049, 50.29292, 45.87027, 42.63018, 39.95224, 38.80347,
    38.15901, 38.0563,
  66.51456, 59.90791, 57.61464, 58.44738, 62.3904, 63.03371, 66.72939,
    69.35304, 75.77998, 78.39835, 68.58653, 63.95237, 70.78558, 70.73927,
    68.36534, 66.1835, 64.32426, 63.26242, 63.73676, 63.2432, 62.7202,
    61.26859, 59.9383, 58.79307, 52.1589, 44.24337, 40.22331, 39.28553,
    38.23899, 38.02334,
  64.91125, 61.94724, 57.64106, 58.73324, 65.60281, 68.47012, 68.65944,
    66.92706, 70.37183, 69.35275, 59.3102, 61.23273, 63.7973, 63.22564,
    60.64481, 60.38786, 59.73927, 57.25844, 57.45063, 58.15379, 58.35842,
    57.40216, 55.92616, 57.83039, 57.39312, 48.7253, 42.04505, 41.38415,
    39.4434, 38.16783,
  70.19398, 69.35551, 69.69067, 72.37937, 75.60075, 74.8857, 77.19713,
    75.89747, 77.37061, 68.98254, 58.40239, 63.06148, 64.52467, 65.59065,
    64.04935, 63.31979, 63.16764, 60.42664, 57.76178, 57.35156, 56.47794,
    55.05785, 54.04552, 54.36851, 55.50557, 54.57926, 48.75156, 43.13465,
    41.04672, 38.91042,
  75.46965, 77.2028, 71.71874, 72.44511, 75.49693, 75.28574, 74.26395,
    76.09195, 80.98473, 72.14986, 58.8508, 64.19929, 65.93971, 67.96163,
    67.52418, 67.1861, 64.81125, 62.82782, 59.74805, 56.51283, 56.21454,
    55.85033, 53.59909, 51.64233, 51.46087, 54.4777, 54.28223, 48.16816,
    44.58585, 41.38755,
  86.58006, 90.23759, 86.1462, 79.99489, 76.97523, 76.03047, 81.88551,
    86.72108, 80.94681, 68.67253, 64.65809, 68.22374, 70.30795, 68.93524,
    65.86289, 65.57517, 64.26189, 62.82639, 61.16457, 58.03984, 57.49844,
    56.20657, 52.24075, 50.01628, 51.18248, 53.4964, 55.5801, 51.54029,
    44.29082, 41.07642,
  95.83875, 94.78203, 83.48343, 77.40009, 76.3495, 76.174, 84.66338,
    84.74379, 73.07624, 65.20995, 68.25743, 70.03402, 69.66871, 66.82285,
    64.48868, 63.35134, 61.85547, 61.11193, 60.24975, 58.53302, 60.24739,
    63.10818, 62.27119, 59.19502, 58.58422, 59.91549, 62.28651, 58.1373,
    45.10635, 38.70855,
  95.35763, 87.6003, 80.14035, 80.4246, 84.27367, 84.52161, 86.23694,
    78.84541, 66.00586, 66.78469, 68.55339, 69.0302, 67.91597, 66.13863,
    65.58386, 63.896, 61.53076, 62.85333, 66.00938, 68.85127, 70.46462,
    69.11379, 64.9033, 62.28544, 61.62729, 62.4173, 62.9452, 64.59501,
    57.40705, 42.62672,
  79.7856, 75.76401, 81.60645, 90.93513, 94.42792, 96.33351, 87.37079,
    69.74047, 61.39735, 62.154, 59.72367, 58.87461, 60.32087, 63.01561,
    66.30329, 68.78821, 70.52997, 72.72615, 71.25916, 67.97832, 66.18161,
    62.63609, 58.57446, 56.19358, 56.49279, 57.13519, 56.28651, 54.05336,
    52.09754, 45.05409,
  80.40018, 83.07077, 85.14417, 85.61212, 89.20976, 95.27397, 91.34602,
    71.57475, 61.43713, 65.69269, 68.54085, 72.03642, 74.60487, 75.32211,
    75.00515, 73.71721, 69.59632, 64.52767, 61.50946, 58.04027, 54.61316,
    52.65774, 51.06731, 49.92416, 49.73685, 50.07961, 48.98944, 45.74913,
    42.3075, 38.62473,
  42.91904, 44.1357, 45.31458, 46.73385, 47.99008, 49.42085, 50.93302,
    52.54615, 54.11284, 55.95846, 58.55074, 59.2174, 56.48892, 57.04771,
    57.11333, 55.69907, 55.05465, 55.03876, 55.07272, 55.98171, 56.1879,
    54.34053, 54.65043, 56.7303, 57.69238, 56.73108, 60.04308, 61.41416,
    47.14188, 41.88303,
  47.43858, 49.53004, 50.28703, 52.82186, 53.79489, 55.03288, 57.11241,
    59.01821, 60.93421, 63.01486, 65.43433, 68.21439, 69.94084, 68.30048,
    66.85004, 67.07552, 65.84548, 66.44459, 67.37875, 68.33888, 68.03768,
    66.81785, 66.2812, 68.37279, 70.69427, 64.87054, 57.40102, 60.4886,
    47.46493, 43.09592,
  51.10638, 53.66103, 55.6731, 57.52666, 58.92596, 60.27116, 61.48384,
    62.7617, 64.04853, 65.228, 66.56418, 68.43855, 70.2791, 72.35167,
    73.28584, 71.07149, 71.8735, 73.91176, 75.68011, 79.10934, 85.0528,
    90.17013, 89.70462, 85.90549, 81.88651, 75.97894, 68.33933, 57.97756,
    46.81281, 43.97453,
  58.61182, 61.33681, 64.26814, 67.04243, 68.89552, 70.87095, 71.60771,
    71.53003, 72.17326, 72.60032, 72.57756, 73.10835, 72.63778, 71.55195,
    74.31534, 75.51411, 72.22694, 70.04355, 74.21303, 79.09686, 86.28227,
    86.72337, 82.23924, 86.92578, 85.35123, 83.48782, 79.42703, 65.18989,
    51.11482, 43.21532,
  68.62782, 70.11713, 73.07021, 75.21511, 76.25491, 76.82763, 77.94911,
    78.74527, 80.66402, 82.01687, 82.23296, 84.75067, 85.84361, 84.68053,
    84.37463, 84.31784, 79.87057, 73.50924, 74.01685, 79.16614, 78.22331,
    69.16335, 70.93195, 77.48293, 83.26199, 83.68694, 80.58332, 85.94633,
    76.61272, 51.05323,
  76.1913, 80.42313, 84.23413, 87.72977, 86.71457, 85.9643, 88.73907,
    89.32015, 88.16151, 89.0053, 92.67491, 101.8147, 110.3488, 107.1952,
    107.4757, 108.7956, 105.0526, 94.0117, 81.84319, 78.67349, 70.18385,
    62.51658, 67.32523, 71.7148, 76.47157, 76.42493, 76.16164, 89.30119,
    80.32136, 46.55054,
  74.54857, 79.37102, 84.08617, 88.80572, 90.54668, 93.42031, 99.69336,
    104.2552, 102.2571, 96.71778, 92.32484, 84.34029, 75.61253, 76.7419,
    78.15971, 80.36749, 80.3217, 75.16538, 68.57368, 68.88385, 65.8931,
    64.63004, 67.67206, 72.45147, 72.73355, 68.05322, 71.56199, 78.42725,
    65.78243, 40.47887,
  74.94423, 80.72279, 86.79261, 92.45195, 95.70976, 103.9278, 107.5256,
    92.05136, 84.35364, 85.58121, 83.37313, 80.78661, 78.61571, 78.53411,
    78.20958, 79.18022, 80.29581, 77.35649, 71.5021, 70.08747, 69.79602,
    71.79434, 75.67307, 76.9746, 72.54681, 71.41659, 77.2328, 74.32584,
    56.64485, 41.58294,
  94.19545, 98.17305, 100.9493, 103.5496, 105.5712, 108.3101, 100.4563,
    100.7311, 104.4651, 105.4794, 105.3171, 104.4347, 104.3548, 109.9361,
    110.8912, 97.43748, 94.47246, 94.45294, 90.14845, 81.76646, 77.93036,
    83.1993, 89.14985, 85.82747, 77.37079, 81.12288, 79.65971, 65.59586,
    43.86688, 41.33387,
  117.9494, 119.9175, 118.3225, 118.3042, 119.9956, 111.5738, 94.33463,
    100.6515, 98.85526, 100.3068, 103.0875, 108.1818, 105.6129, 101.4983,
    97.37476, 101.5504, 101.314, 96.98113, 91.29884, 89.08173, 90.44286,
    85.71748, 79.24623, 70.96359, 75.14261, 82.20291, 71.63685, 50.3975,
    40.84204, 39.25851,
  118.8089, 118.3025, 119.9253, 119.6634, 120.8208, 119.1359, 108.4212,
    108.1725, 107.6372, 101.4625, 88.31862, 71.70921, 69.23013, 69.93546,
    70.74635, 72.49263, 74.76856, 75.25013, 75.08678, 77.56599, 85.37749,
    79.9789, 66.56885, 63.77787, 67.44289, 63.50151, 49.8001, 41.86589,
    41.38256, 39.41605,
  125.0354, 121.6841, 124.5227, 124.725, 123.4583, 119.3941, 112.6693,
    103.3103, 94.90219, 85.49319, 79.68928, 75.97871, 78.17503, 78.06973,
    73.68073, 71.3156, 68.78048, 68.00217, 67.82362, 71.20386, 78.194,
    75.13044, 65.27309, 72.82477, 74.09818, 58.53849, 42.84929, 45.89753,
    42.72699, 40.53482,
  126.9452, 127.6009, 129.5208, 130.3757, 129.3183, 126.2041, 120.286,
    117.4114, 118.7454, 112.6367, 105.4639, 97.99032, 103.0698, 103.9199,
    92.28992, 77.71201, 77.01966, 74.17589, 71.92484, 74.27831, 75.04088,
    68.31142, 62.21841, 58.96523, 58.04305, 51.36654, 43.97944, 44.97618,
    44.35223, 41.62831,
  115.9385, 117.3966, 118.3222, 118.5248, 118.7941, 119.9236, 121.3217,
    121.8007, 119.8345, 119.783, 120.2769, 118.9175, 119.7355, 119.9086,
    113.7976, 95.16417, 87.2419, 89.16379, 89.55257, 80.61162, 69.54179,
    62.04871, 56.91379, 49.49042, 45.63886, 44.73026, 42.44275, 41.48481,
    41.87302, 41.002,
  111.5297, 109.5025, 112.9665, 114.6978, 116.3711, 119.0755, 121.3192,
    121.2829, 113.4965, 111.7964, 105.7425, 100.2309, 101.5743, 104.4554,
    103.2511, 99.0571, 89.37852, 84.27685, 81.8943, 73.90005, 59.05378,
    56.90024, 50.16057, 47.42928, 46.47022, 44.81671, 42.87854, 41.45604,
    40.51845, 39.94345,
  110.2879, 114.241, 115.242, 114.4296, 113.1304, 114.7138, 116.9326,
    109.8402, 99.94894, 94.38913, 92.12187, 86.36108, 82.87428, 88.77438,
    85.53671, 82.32968, 81.93265, 73.91685, 70.47099, 63.08739, 51.67194,
    52.4952, 47.88784, 46.2964, 45.89571, 44.38465, 42.50739, 41.52583,
    40.66874, 39.94464,
  94.08183, 92.95572, 94.5622, 96.85043, 98.69672, 101.4859, 104.3213,
    106.7329, 105.5037, 99.24907, 91.27924, 97.87218, 103.7883, 94.73461,
    88.07736, 81.02112, 75.14813, 71.15757, 69.97514, 63.92706, 51.97383,
    52.8469, 48.64753, 46.1947, 44.97535, 44.20918, 41.79808, 40.135,
    40.0389, 39.76154,
  85.48252, 85.90352, 84.09086, 86.00885, 88.25538, 91.8654, 95.21646,
    99.19134, 102.0138, 102.2881, 109.5901, 114.7948, 110.5087, 109.2861,
    103.0242, 93.37435, 83.21347, 79.96413, 79.81503, 69.4372, 53.92794,
    52.06176, 48.68462, 46.89648, 43.8368, 42.64714, 41.64371, 39.677,
    39.57895, 39.42606,
  93.32761, 84.67755, 75.08685, 70.9966, 74.41699, 76.75385, 80.22557,
    83.3635, 84.79094, 87.77457, 92.45939, 90.35415, 83.8002, 88.1556,
    90.37427, 92.25641, 98.48926, 102.9215, 98.46882, 84.34866, 64.63074,
    55.30233, 50.48381, 47.41941, 44.0418, 42.13068, 41.30792, 40.05164,
    39.57792, 39.44454,
  87.41063, 80.7637, 73.16797, 68.78448, 71.57745, 73.14273, 74.76279,
    75.95037, 78.14404, 82.74669, 81.57743, 71.61606, 71.86822, 71.67529,
    70.54824, 70.03873, 74.54388, 81.14834, 83.32391, 80.91402, 72.27019,
    62.06322, 54.3144, 50.31842, 46.77346, 43.11985, 41.63377, 40.30009,
    39.59865, 39.46889,
  84.00468, 78.40645, 70.63605, 66.373, 66.80838, 66.90364, 67.34354,
    68.42522, 70.94235, 73.0893, 68.07525, 61.85293, 66.27226, 65.64486,
    63.19748, 61.46943, 62.63663, 64.65738, 66.83573, 66.93832, 66.44084,
    66.15981, 61.35727, 54.95456, 49.46264, 44.50528, 41.63808, 40.45401,
    39.61198, 39.47664,
  86.89655, 79.93874, 72.00845, 68.1823, 67.36752, 64.72006, 65.4917,
    66.1599, 70.04513, 69.95937, 62.17759, 58.42797, 61.16642, 60.92682,
    59.58406, 58.98765, 58.25168, 58.63191, 60.30629, 60.99971, 60.90742,
    60.64248, 61.4364, 61.12365, 55.22352, 46.54149, 42.56536, 41.40613,
    39.89331, 39.46864,
  90.59025, 87.40149, 77.83279, 74.94498, 77.93441, 77.83622, 76.14276,
    73.03236, 73.16459, 70.15415, 62.94635, 64.25191, 65.4151, 65.21895,
    63.40429, 63.11609, 61.73349, 58.64055, 57.69201, 57.47149, 57.05878,
    56.65946, 56.31494, 58.91697, 60.09751, 52.59315, 45.50471, 43.77596,
    41.54792, 39.66905,
  96.58451, 94.61412, 90.16965, 90.12189, 89.90421, 88.84589, 90.01026,
    89.04581, 90.02088, 81.72861, 74.29511, 77.82361, 79.29499, 79.61209,
    76.5565, 73.87953, 71.27332, 66.57475, 62.13032, 60.1465, 58.14829,
    56.74063, 55.95168, 56.00108, 58.05366, 58.78095, 53.5363, 46.70578,
    44.03863, 40.84145,
  96.82596, 93.35567, 85.81961, 84.00658, 85.35051, 84.14146, 84.85951,
    88.86241, 92.74331, 84.28782, 76.1978, 79.34259, 80.63656, 81.35679,
    79.69604, 77.92252, 73.98195, 70.62611, 67.46992, 63.82507, 61.58429,
    59.04866, 55.91225, 54.02845, 54.93943, 58.0048, 58.75457, 51.43557,
    46.49908, 42.91302,
  102.8571, 100.6719, 94.90403, 88.10072, 85.47314, 84.27525, 88.83573,
    93.5688, 91.30643, 83.90012, 83.29361, 84.25438, 84.54337, 82.61903,
    79.60775, 78.18337, 75.97084, 73.74228, 72.63656, 70.33563, 68.70147,
    66.58498, 62.15338, 58.74902, 58.70346, 60.17574, 61.49164, 54.28418,
    44.87598, 41.76068,
  102.1931, 97.79417, 90.08108, 86.32349, 84.28143, 82.01665, 86.79613,
    88.26157, 85.06348, 82.94772, 85.28553, 85.77438, 84.53944, 82.70294,
    80.14385, 77.33778, 74.66975, 73.30095, 72.92067, 71.71363, 71.51475,
    72.49052, 71.27313, 67.77798, 67.05119, 69.22964, 72.16649, 65.30567,
    48.88943, 40.28177,
  100.8258, 96.37379, 94.68056, 94.34825, 95.38737, 92.01106, 89.4341,
    83.99107, 77.10954, 77.51831, 77.57175, 78.06429, 77.97874, 77.19444,
    76.21577, 73.0677, 68.86862, 67.24548, 67.84416, 68.07198, 65.60009,
    62.18063, 59.3959, 58.46349, 60.06669, 62.69739, 64.82934, 67.00305,
    60.33557, 44.61023,
  87.01698, 86.50083, 89.65478, 93.0881, 96.29102, 97.22256, 87.61295,
    74.20096, 68.60211, 68.45834, 66.23576, 65.3886, 65.39227, 65.09933,
    64.58051, 63.20369, 60.73914, 58.53623, 55.94948, 52.91886, 51.5647,
    50.59882, 48.60893, 47.36525, 48.75994, 50.30732, 50.22704, 48.97953,
    49.45755, 45.27468,
  71.04898, 72.35345, 70.95154, 69.79617, 73.32137, 79.30807, 78.23711,
    64.96202, 58.64711, 62.02996, 63.87118, 65.2321, 65.28069, 62.87937,
    59.77547, 56.89632, 51.83823, 46.98214, 46.20691, 45.40633, 43.78175,
    44.01532, 44.05745, 44.00212, 44.44481, 45.59248, 45.70294, 43.63781,
    41.43102, 39.49089,
  54.28894, 54.71279, 55.04905, 55.48284, 55.56351, 55.83839, 56.3041,
    56.84197, 57.42741, 58.34319, 59.7532, 59.61835, 57.01146, 57.02288,
    56.88595, 55.93689, 55.63531, 55.87471, 56.1236, 56.75953, 56.54434,
    54.83759, 54.97327, 56.65533, 57.60461, 56.7239, 58.51018, 59.89629,
    49.69228, 45.85414,
  59.80487, 60.26855, 59.78956, 60.6109, 60.2672, 60.18555, 60.83678,
    61.55429, 62.47597, 63.62217, 65.01859, 66.70807, 67.70613, 66.26414,
    65.20456, 65.57862, 65.12399, 65.96465, 66.92702, 67.61758, 67.10225,
    65.80503, 64.89371, 66.50692, 68.20602, 62.64582, 55.83315, 58.71489,
    50.17384, 46.73522,
  61.97742, 62.2286, 62.25077, 62.24531, 62.07377, 62.06284, 62.02273,
    62.17552, 62.53355, 63.04804, 63.75824, 65.07496, 66.616, 68.17233,
    69.07788, 68.16355, 69.39044, 71.66402, 73.83159, 76.97835, 82.03449,
    86.1474, 84.92766, 80.62769, 76.9027, 71.97062, 65.11543, 57.48875,
    49.52142, 47.39325,
  67.54889, 67.77106, 68.26364, 68.78646, 69.08838, 69.60178, 69.3121,
    68.52464, 68.541, 68.42969, 67.91458, 68.07296, 67.59132, 66.74515,
    68.79832, 70.20879, 68.47057, 67.52296, 71.28765, 75.6283, 82.30202,
    83.17171, 78.04774, 80.81894, 78.48428, 77.01524, 75.05328, 63.99162,
    52.81107, 46.82898,
  72.82706, 72.35345, 73.10646, 73.38659, 73.2589, 73.06662, 73.40707,
    73.40996, 74.62454, 75.43223, 75.46841, 77.70842, 78.87762, 77.93817,
    77.7721, 78.09981, 75.01971, 70.6534, 70.98047, 75.33028, 75.06258,
    66.92916, 68.23167, 72.96013, 77.2457, 77.8997, 75.83603, 81.29164,
    75.40509, 53.90028,
  76.70645, 78.8838, 80.52666, 82.03763, 80.96001, 80.60666, 82.8455,
    82.87178, 81.33174, 80.87181, 82.72798, 89.85918, 97.53122, 95.49925,
    96.02652, 97.00117, 94.71104, 87.3644, 77.82261, 74.88013, 67.93605,
    61.53326, 65.30025, 68.41057, 72.31706, 73.03421, 73.45167, 85.12036,
    79.25288, 50.02213,
  81.10104, 84.05223, 86.32896, 88.40805, 88.88721, 91.16616, 96.57312,
    100.0119, 97.98391, 92.24358, 86.95355, 77.98174, 68.95634, 69.91211,
    71.04543, 73.3471, 74.49863, 72.12357, 67.61752, 67.28835, 64.2489,
    63.02974, 65.34656, 68.88033, 69.37347, 66.27975, 69.08418, 76.08548,
    66.74593, 44.53477,
  83.24435, 85.96384, 88.81133, 91.45151, 92.51848, 98.16429, 100.5682,
    85.94922, 78.33649, 78.71061, 75.826, 72.7186, 70.70871, 70.7766,
    70.67471, 71.82019, 74.41601, 73.7094, 69.64548, 68.18781, 67.31382,
    68.46938, 71.19437, 72.5639, 70.11014, 69.26897, 73.96582, 72.35062,
    57.62709, 45.36639,
  88.94004, 88.82502, 88.49796, 89.16959, 89.58717, 90.17098, 81.23119,
    80.16253, 82.38918, 83.23327, 83.57465, 83.10123, 83.43355, 88.22009,
    90.55632, 82.99784, 82.57857, 84.0472, 81.92706, 76.2739, 72.58841,
    75.71594, 79.72585, 78.03568, 73.18393, 76.7741, 76.37198, 65.55987,
    47.21242, 45.51737,
  111.4215, 109.8456, 99.52527, 97.55241, 96.87692, 89.47563, 73.54735,
    77.78145, 76.02613, 77.00037, 78.48582, 82.11215, 80.87186, 79.34769,
    78.09545, 82.28693, 83.7757, 82.41919, 80.30988, 79.43093, 80.21558,
    76.58724, 72.18604, 66.6246, 70.50919, 77.93813, 70.79201, 52.42103,
    45.16528, 43.97577,
  121.0246, 119.8401, 119.5196, 114.8461, 113.7266, 101.5242, 91.57507,
    89.6236, 88.72053, 85.52127, 75.63543, 63.52784, 62.10373, 62.53492,
    63.20307, 64.76558, 66.87914, 68.29932, 69.15822, 71.34666, 77.24696,
    73.9781, 64.73279, 62.8546, 66.22549, 64.50018, 52.66069, 45.66361,
    45.51618, 44.09585,
  127.841, 124.7378, 125.4115, 124.5119, 121.6561, 113.8549, 104.0208,
    93.9109, 86.93129, 80.69206, 75.44882, 71.74539, 72.99913, 71.79512,
    66.85006, 65.43275, 64.32628, 64.3616, 64.65857, 67.41377, 72.82909,
    71.42535, 64.16566, 70.17234, 72.91157, 60.21645, 46.58819, 49.12895,
    46.51439, 44.90229,
  123.6173, 124.5478, 125.3681, 125.6946, 125.2901, 122.6459, 116.1447,
    107.7777, 111.4826, 101.4471, 95.14923, 89.77341, 93.40244, 93.50446,
    82.80846, 70.10761, 70.70721, 69.5994, 68.04551, 69.33181, 70.49247,
    66.75446, 62.48961, 59.17743, 58.91624, 54.20422, 47.74673, 48.53792,
    47.92865, 45.80592,
  101.5797, 102.7743, 98.07273, 97.84919, 99.1772, 107.4301, 115.9366,
    115.1879, 103.2711, 106.1114, 111.4771, 105.6934, 106.5072, 105.9702,
    96.5405, 83.54468, 77.45887, 80.30867, 81.38342, 75.01595, 67.40542,
    62.0711, 57.37882, 51.47913, 48.19902, 48.10262, 46.53076, 45.72389,
    45.93887, 45.29533,
  85.017, 81.52592, 82.24414, 82.17888, 82.88587, 84.73729, 88.99216,
    88.45689, 84.01137, 84.88876, 81.63516, 79.39482, 81.30829, 85.23973,
    86.36035, 85.31783, 79.47617, 75.10627, 73.01814, 68.67464, 59.14169,
    57.24182, 51.65222, 49.25581, 48.95758, 48.04995, 46.79375, 45.63908,
    44.86309, 44.42248,
  86.96624, 89.4361, 89.98871, 89.30443, 87.79908, 89.41341, 91.02182,
    85.82246, 81.21555, 76.81447, 76.04269, 72.7339, 70.76328, 74.46086,
    72.4124, 71.20937, 72.12925, 67.31854, 64.45781, 59.89052, 52.953,
    53.15068, 49.65081, 48.71855, 48.61236, 47.85988, 46.56418, 45.63217,
    44.92834, 44.42929,
  77.01698, 76.25975, 77.4837, 79.48874, 81.25883, 83.01342, 85.30305,
    88.04109, 86.62576, 83.2875, 78.94931, 83.5248, 87.83068, 82.38071,
    76.22715, 71.29633, 67.60428, 65.30649, 64.33102, 60.57169, 53.18902,
    53.55683, 50.4276, 48.84272, 48.20677, 47.69502, 46.012, 44.69372,
    44.55289, 44.32837,
  69.35461, 69.25251, 68.14317, 70.06906, 72.17778, 74.79459, 77.06636,
    79.57823, 81.6348, 81.85062, 86.96729, 91.15257, 90.39528, 91.14526,
    87.04944, 81.62861, 76.03449, 74.118, 73.02216, 65.4564, 54.95368,
    53.10115, 50.73016, 49.5542, 47.4991, 46.62361, 45.86089, 44.34052,
    44.21737, 44.06478,
  75.29588, 69.10431, 61.81742, 58.28914, 60.59148, 61.52814, 63.47018,
    65.50865, 66.36502, 68.9395, 72.94452, 72.0979, 68.82384, 72.35699,
    74.78675, 77.43856, 83.44395, 88.12794, 85.87574, 77.07375, 63.68251,
    55.85692, 51.86561, 49.93811, 47.69455, 46.33416, 45.6106, 44.55676,
    44.18655, 44.08438,
  72.38545, 66.85043, 59.57392, 55.11013, 56.41571, 57.21991, 58.50858,
    59.86676, 62.13958, 66.25232, 66.79912, 61.23311, 61.80579, 61.27678,
    60.75885, 61.5323, 65.52112, 71.14249, 73.39649, 72.56061, 67.34533,
    60.15263, 54.56838, 51.98766, 49.72519, 47.11099, 45.82345, 44.69049,
    44.18341, 44.10759,
  73.75481, 69.10278, 61.33019, 56.93462, 56.76187, 56.76013, 57.45841,
    58.52767, 60.63298, 62.85398, 60.37844, 56.69392, 59.66261, 59.37536,
    58.15818, 57.63875, 58.98623, 60.7886, 62.51739, 62.1883, 61.70461,
    61.74164, 59.03004, 55.18481, 51.55812, 48.03256, 45.85966, 44.74928,
    44.16409, 44.1148,
  80.97882, 77.36308, 69.60096, 65.8844, 64.99039, 62.52753, 62.0915,
    61.67672, 63.70726, 63.89794, 59.18822, 56.66024, 58.27904, 58.14364,
    57.53107, 57.47264, 57.22821, 57.64231, 58.85713, 59.14303, 58.90507,
    58.81275, 59.5848, 59.42897, 55.23936, 49.34281, 46.54333, 45.46,
    44.36382, 44.06366,
  86.6378, 86.43712, 78.20319, 75.23822, 76.65411, 76.03271, 73.76345,
    70.53687, 70.25462, 68.09107, 63.26536, 63.54142, 63.83903, 63.43668,
    61.77465, 61.37307, 60.67904, 58.65368, 57.97148, 57.61322, 56.91838,
    56.63211, 56.54955, 57.94832, 58.45644, 53.4835, 48.75418, 47.14028,
    45.49624, 44.2316,
  88.9968, 88.39973, 83.52934, 81.51766, 81.35978, 80.20634, 80.63938,
    80.27137, 81.7003, 77.0014, 72.00172, 73.86075, 74.80368, 74.63585,
    72.19135, 70.12527, 68.44894, 65.55471, 62.2953, 60.35467, 58.39837,
    57.15775, 56.41816, 56.22848, 57.63398, 58.1608, 54.36343, 49.36663,
    47.47722, 45.13888,
  90.26974, 85.5631, 79.05812, 76.23746, 76.11897, 75.55886, 76.49023,
    79.58903, 83.26141, 78.43557, 72.86697, 74.62488, 75.67743, 75.92255,
    74.64493, 73.6318, 71.64005, 69.74393, 66.82584, 63.71288, 61.65823,
    59.68015, 57.02941, 55.46968, 56.31504, 58.24069, 57.97938, 52.46798,
    49.14293, 46.60202,
  91.53128, 87.7301, 82.00488, 76.1125, 73.64153, 72.70709, 76.07995,
    79.90939, 79.28416, 74.43298, 74.10886, 74.96581, 75.73847, 74.97713,
    73.25515, 72.98208, 72.77402, 72.04163, 70.43237, 68.14111, 66.86926,
    65.3243, 61.58869, 59.02168, 59.04129, 58.93471, 58.77393, 54.18108,
    47.95826, 45.7122,
  87.33543, 83.14329, 76.85813, 72.20203, 69.47379, 66.85044, 69.80907,
    70.88244, 69.00792, 67.66942, 69.69057, 71.10114, 71.82667, 71.80569,
    71.08346, 70.70526, 70.81065, 71.10933, 70.33858, 69.0345, 68.91475,
    69.48628, 68.3112, 65.85687, 65.04295, 64.78442, 65.12086, 60.88687,
    50.31874, 44.68408,
  79.62853, 77.71188, 74.63054, 73.40224, 72.9371, 69.9785, 67.84401,
    64.37047, 60.64122, 61.53982, 62.67714, 64.38132, 66.04195, 66.92843,
    67.46126, 66.93626, 65.79485, 65.59035, 65.74284, 65.52563, 64.06317,
    62.05026, 59.88943, 59.2705, 60.15823, 60.93991, 61.34049, 62.16942,
    57.5822, 47.52363,
  65.10868, 64.78174, 66.09305, 67.91373, 70.73208, 72.80971, 68.13458,
    59.74237, 57.29798, 58.50204, 58.20927, 58.35277, 59.21059, 59.94601,
    60.26251, 60.00462, 59.04741, 58.01659, 56.16578, 54.11706, 53.45872,
    52.81998, 51.60667, 50.95547, 51.96233, 52.95508, 52.70588, 51.28109,
    50.97184, 48.03087,
  56.39863, 56.78394, 56.37023, 56.10518, 58.95982, 64.11044, 64.80592,
    56.91173, 53.29163, 55.95065, 57.64573, 58.94119, 59.30923, 58.04233,
    56.38453, 55.0867, 52.13766, 49.34392, 49.03424, 48.38351, 47.38562,
    47.63671, 47.8511, 47.96077, 48.32611, 49.17282, 49.07824, 47.32653,
    45.62265, 44.12301,
  51.22165, 51.38177, 51.4487, 51.57752, 51.52929, 51.6279, 51.80299,
    52.06017, 52.3882, 52.9255, 53.81587, 53.30859, 50.98837, 51.279,
    51.34378, 50.81386, 50.88095, 51.31651, 51.82601, 52.71553, 53.15718,
    52.33881, 52.97378, 54.84925, 56.00629, 55.26917, 56.21809, 57.11674,
    49.3357, 46.44032,
  56.58526, 56.95422, 56.4003, 56.94422, 56.60057, 56.38659, 56.69308,
    56.97403, 57.32557, 57.72565, 58.27704, 58.90445, 59.13306, 57.78643,
    56.77237, 57.0971, 56.54115, 57.08443, 57.91906, 58.68996, 58.7965,
    58.79959, 59.70851, 62.98838, 65.86687, 61.00326, 53.66557, 56.74278,
    49.63497, 47.16008,
  58.3824, 58.85216, 59.05956, 59.25764, 59.41662, 59.66423, 59.93191,
    60.40988, 60.95825, 61.40562, 61.9178, 62.77714, 63.70697, 64.76593,
    65.33522, 64.46344, 65.19061, 66.66785, 68.11603, 70.55777, 75.12209,
    79.69423, 79.75506, 76.50938, 73.82682, 68.74195, 62.63668, 55.95093,
    49.7173, 47.99359,
  61.84879, 62.30759, 63.06743, 63.89421, 64.4302, 65.09777, 65.14315,
    64.69742, 64.91681, 65.15872, 65.11405, 65.55893, 65.63682, 65.32181,
    67.39897, 68.75323, 67.41708, 66.55227, 69.76059, 73.75443, 79.7039,
    79.72429, 73.78833, 75.82799, 73.25392, 71.0867, 69.24996, 59.82764,
    51.05753, 47.1324,
  66.79333, 66.73175, 67.68066, 68.33153, 68.62064, 68.71992, 69.05347,
    69.02607, 69.84756, 70.11441, 69.93259, 71.34192, 72.31977, 72.18396,
    72.83401, 73.8303, 72.1854, 69.4181, 71.01346, 75.82982, 75.86976,
    67.40225, 67.12254, 71.39391, 74.46237, 74.48148, 73.00598, 77.86829,
    72.9969, 54.63934,
  72.46329, 74.7354, 76.62556, 78.51196, 78.36372, 78.85303, 81.31159,
    82.02847, 81.92087, 82.82892, 85.47227, 92.5659, 99.91632, 97.66057,
    98.47557, 99.69695, 95.97779, 87.87173, 78.78204, 75.87898, 69.35658,
    62.63735, 66.5955, 69.8576, 73.80003, 75.05259, 76.47878, 86.68813,
    80.18221, 51.16137,
  74.48557, 77.14164, 79.42293, 81.69077, 82.81362, 85.97062, 92.0946,
    96.91663, 96.25585, 91.63039, 87.53934, 79.76476, 71.39105, 72.52777,
    73.61919, 75.1228, 75.59239, 71.95715, 66.83101, 66.0118, 63.03658,
    62.01435, 64.609, 68.0724, 69.12115, 67.55995, 71.62447, 77.56082,
    66.71358, 45.34274,
  74.08994, 76.52699, 78.9711, 81.58623, 83.04587, 88.33458, 91.12547,
    78.12555, 70.98862, 71.04232, 68.34145, 65.5006, 63.95504, 64.70709,
    65.6749, 67.70813, 69.97794, 69.13206, 65.62593, 64.60438, 63.9802,
    65.16008, 67.92644, 69.92444, 68.92081, 69.44984, 74.5906, 72.55965,
    58.36142, 45.73102,
  80.11744, 81.65767, 82.75171, 83.97339, 85.51614, 87.03567, 78.92077,
    77.45934, 79.57916, 79.70212, 79.361, 78.51533, 79.15501, 83.44147,
    85.55463, 80.05376, 80.46378, 81.81602, 79.7339, 74.20077, 71.20337,
    74.05247, 77.4214, 76.23377, 72.93043, 77.58034, 78.00294, 66.79021,
    47.78628, 46.30591,
  93.97508, 96.18466, 90.34413, 90.02219, 92.00915, 87.22553, 72.34506,
    77.53516, 77.06898, 79.01625, 80.71835, 84.21741, 83.35464, 81.63821,
    79.79276, 82.51473, 83.10014, 81.48882, 79.37067, 77.90121, 78.31334,
    75.52052, 72.12602, 68.09302, 72.52064, 79.60073, 72.33774, 53.56564,
    45.78413, 45.00639,
  107.3587, 106.7194, 107.1208, 99.49337, 99.94562, 90.26625, 81.22845,
    82.56784, 83.66798, 81.39703, 73.30688, 63.65755, 62.87931, 63.65693,
    63.93527, 65.24572, 66.74429, 67.33018, 67.66856, 69.15664, 74.00526,
    71.4592, 64.01735, 62.94722, 67.19163, 66.01632, 54.18, 46.16083,
    46.4654, 45.03767,
  114.4357, 111.2835, 112.9794, 112.1229, 109.4776, 96.15811, 90.4931,
    82.36919, 76.23235, 72.70399, 68.72125, 66.5144, 68.60553, 67.98576,
    64.74493, 64.3768, 63.64844, 63.79554, 64.03074, 66.32234, 71.26828,
    70.75784, 64.82373, 70.59868, 72.66351, 60.37369, 47.08802, 49.58664,
    47.23993, 45.8702,
  116.2606, 116.8495, 117.7225, 117.0828, 115.0141, 111.407, 105.0822,
    96.32287, 100.8911, 90.25722, 84.70197, 79.91779, 83.95325, 85.01699,
    77.74236, 67.27892, 67.76826, 67.18618, 66.42905, 68.22333, 70.1849,
    68.24045, 65.00735, 62.02149, 60.46985, 55.00662, 48.70663, 49.60847,
    48.70433, 46.71384,
  106.4014, 107.1204, 106.8689, 105.5384, 104.8319, 105.2334, 105.6537,
    105.2003, 103.1083, 102.8279, 102.8319, 101.6445, 101.1442, 101.3382,
    93.73428, 80.0356, 76.11245, 78.55962, 79.93814, 74.08808, 66.90669,
    62.56697, 58.85611, 52.74274, 49.36623, 48.92227, 47.46534, 46.79022,
    46.85526, 46.20528,
  82.20367, 79.48736, 81.70287, 82.28407, 83.83124, 86.85326, 92.22989,
    91.54074, 87.26024, 87.34883, 84.06204, 80.33943, 82.21659, 85.23868,
    85.22069, 84.52692, 77.57358, 74.47795, 72.37598, 67.83662, 58.64371,
    56.53475, 51.7411, 49.53482, 49.39019, 48.71125, 47.40472, 46.41581,
    45.74943, 45.38669,
  79.16004, 81.24644, 81.89403, 81.45373, 80.40825, 81.66175, 83.71764,
    80.61102, 76.09074, 73.20323, 72.64929, 70.49848, 69.66681, 73.09954,
    71.14661, 69.51225, 69.96872, 65.57881, 63.09145, 58.82681, 52.4066,
    52.56979, 49.68032, 48.8136, 48.90399, 48.41422, 47.27275, 46.54784,
    45.85872, 45.36877,
  72.87865, 72.02315, 72.63559, 73.83071, 74.89537, 75.85766, 77.15987,
    78.99231, 78.05895, 75.30029, 71.3469, 75.10006, 79.46465, 75.66351,
    70.59045, 67.40489, 64.45094, 62.46001, 61.95108, 59.23251, 52.84737,
    52.90372, 50.09772, 48.93182, 48.63786, 48.3068, 46.91796, 45.79985,
    45.51733, 45.31715,
  69.47254, 70.06017, 69.19295, 70.60617, 71.93852, 73.58627, 75.02267,
    76.89215, 78.47846, 77.50296, 80.54701, 83.40083, 82.29778, 81.52724,
    76.53166, 72.38903, 67.48911, 65.97542, 66.30782, 61.3819, 53.16515,
    52.19131, 50.27702, 49.48818, 48.15007, 47.43479, 46.73737, 45.41496,
    45.24924, 45.09326,
  77.63756, 73.01028, 66.31149, 63.32178, 65.66797, 66.46935, 68.07451,
    69.96992, 70.56284, 72.44533, 75.53252, 74.78017, 71.16191, 72.85929,
    72.94041, 74.5133, 78.95815, 82.22623, 80.24372, 72.25903, 60.47786,
    53.69422, 50.6959, 49.73542, 48.23632, 47.20367, 46.53986, 45.60045,
    45.19799, 45.08075,
  73.83295, 69.59095, 62.94386, 59.24751, 60.90295, 61.82372, 63.0842,
    64.42526, 66.44428, 69.71747, 70.09786, 65.48625, 65.66008, 64.66068,
    63.46126, 63.77151, 66.52061, 70.42881, 71.32874, 69.7863, 64.11269,
    57.55032, 53.13055, 51.5569, 49.88739, 47.89889, 46.80828, 45.71917,
    45.1826, 45.11693,
  70.65239, 67.02185, 60.09759, 56.62901, 57.29949, 57.74076, 58.6221,
    59.81859, 61.73805, 63.71857, 61.64631, 58.4351, 60.8952, 60.56744,
    59.0388, 58.13151, 58.87616, 59.92964, 60.81898, 60.119, 59.54331,
    59.158, 56.57154, 53.84626, 51.07624, 48.48822, 46.74489, 45.76033,
    45.17549, 45.10463,
  72.37152, 69.03355, 62.29288, 59.14896, 59.32719, 58.1599, 58.57762,
    58.8805, 61.04063, 61.7259, 58.14109, 56.04514, 57.57708, 57.6687,
    57.09121, 57.08499, 57.08154, 57.57639, 58.40224, 58.84644, 58.84238,
    58.41307, 58.29454, 56.87023, 53.24615, 49.28446, 47.2645, 46.23439,
    45.30062, 45.07729,
  77.45734, 76.30834, 68.58191, 65.78302, 67.15404, 66.98584, 65.63644,
    63.50779, 63.82388, 62.64581, 58.81665, 58.88395, 59.18218, 59.1746,
    58.38924, 58.70577, 58.73339, 57.62704, 57.06477, 56.77773, 56.47524,
    56.14793, 55.44635, 55.42389, 55.48784, 52.25191, 48.77196, 47.58092,
    46.18442, 45.18546,
  81.80028, 81.44046, 76.62318, 74.54124, 74.41966, 72.92799, 73.00658,
    72.88428, 74.58237, 71.7497, 67.83482, 69.01883, 69.38715, 69.1088,
    67.39159, 66.47358, 65.50262, 63.29447, 60.33362, 58.51756, 57.06275,
    56.44814, 55.7608, 54.92435, 55.75236, 56.07808, 53.01818, 49.25703,
    47.75497, 45.95544,
  83.01201, 79.74673, 73.87041, 71.44002, 71.45533, 70.72033, 71.41589,
    73.92403, 77.0029, 73.34557, 68.86304, 70.59705, 71.53588, 71.47891,
    69.85884, 69.55255, 68.25819, 66.65016, 64.04864, 61.44175, 59.61299,
    58.05737, 56.05685, 54.76934, 55.60467, 56.86411, 56.28762, 52.24671,
    49.47377, 47.33791,
  85.23393, 83.01814, 77.65895, 72.8729, 71.60661, 71.16582, 74.06841,
    77.39613, 76.83417, 72.00252, 71.19302, 72.25167, 73.09402, 71.65724,
    69.20556, 68.96817, 68.60437, 67.38864, 65.76641, 63.8067, 62.11758,
    60.367, 57.66941, 56.16198, 56.60102, 56.3315, 56.17503, 53.13869,
    48.56968, 46.63262,
  83.84601, 81.09093, 76.29836, 72.72038, 71.19576, 69.76652, 72.79215,
    74.28276, 72.91136, 71.01942, 72.02025, 73.20457, 73.84167, 72.93133,
    71.26644, 70.71458, 70.15287, 69.19666, 68.05185, 67.00006, 66.45531,
    66.3298, 65.11857, 63.1657, 62.35896, 61.36517, 61.01896, 57.69815,
    49.71652, 45.60347,
  79.21767, 77.51566, 74.97814, 74.5056, 74.66579, 72.93079, 71.86396,
    69.81695, 67.08419, 67.61007, 68.54185, 70.19039, 71.69086, 72.07761,
    71.71267, 70.74861, 69.19389, 68.37625, 68.05846, 67.69322, 65.8251,
    63.18919, 60.95546, 60.0859, 60.36583, 60.22478, 59.81248, 60.13233,
    56.13702, 47.77029,
  67.22279, 67.13567, 68.47803, 70.15178, 72.44424, 73.7545, 69.55634,
    62.88175, 60.84475, 61.2644, 60.75023, 61.13922, 62.44849, 63.62378,
    64.09942, 63.58032, 62.17141, 60.82466, 58.64688, 56.45105, 55.45435,
    54.47408, 53.15298, 52.37428, 53.03996, 53.6729, 53.16554, 51.6871,
    51.1034, 48.43296,
  59.91811, 60.33349, 60.53625, 60.63823, 62.85806, 66.94293, 67.06504,
    60.40639, 57.35505, 59.36685, 60.38741, 61.37681, 61.89212, 61.22879,
    59.75215, 58.17216, 55.11753, 52.36892, 51.60215, 50.5843, 49.54234,
    49.66363, 49.88103, 49.86872, 50.06289, 50.61447, 50.11966, 48.22756,
    46.58328, 45.177,
  50.38474, 50.44233, 50.57504, 50.65535, 50.72771, 50.92733, 51.21397,
    51.59298, 52.02122, 52.56239, 53.36643, 53.10653, 51.45378, 51.75087,
    51.84401, 51.46066, 51.64116, 51.9904, 52.38403, 53.18802, 53.60745,
    53.09743, 53.62745, 55.20206, 56.75537, 56.82904, 57.85457, 58.95887,
    53.50496, 51.34984,
  51.59143, 51.70158, 51.40554, 51.84252, 51.6816, 51.68415, 52.09848,
    52.48344, 52.93296, 53.39291, 53.90916, 54.43758, 54.61762, 53.67041,
    53.10895, 53.67675, 53.5024, 54.3216, 55.34775, 56.2777, 56.63955,
    57.14567, 58.77546, 62.69041, 66.20763, 62.40443, 56.66015, 59.26163,
    53.84993, 51.87329,
  51.68951, 51.73622, 51.84373, 51.95429, 52.05205, 52.26874, 52.53626,
    52.90847, 53.36835, 53.84666, 54.36607, 55.18657, 56.1479, 57.33995,
    58.28563, 58.23573, 59.64135, 61.64317, 63.48428, 66.2482, 70.95833,
    76.17965, 77.54543, 75.63374, 73.75592, 68.7392, 63.91316, 58.639,
    54.01777, 52.64908,
  54.52131, 55.00802, 55.75413, 56.58022, 57.26125, 58.09467, 58.34887,
    58.29288, 58.7073, 59.31442, 59.90567, 61.00511, 61.92835, 62.5303,
    65.14069, 67.32247, 67.18182, 67.29062, 70.66164, 74.90671, 80.92176,
    80.75966, 74.5912, 75.42216, 72.34235, 70.41505, 68.78283, 61.24345,
    54.2003, 51.75219,
  57.62431, 57.37096, 58.15771, 58.69515, 58.99115, 59.13924, 59.5101,
    59.72101, 60.45214, 60.95301, 61.07267, 62.66423, 64.28929, 65.75539,
    67.73975, 70.09772, 70.19627, 69.26721, 72.0015, 76.82923, 76.65296,
    68.71623, 67.38393, 71.06918, 73.16051, 72.7012, 72.01521, 77.3205,
    74.40009, 58.85754,
  59.44811, 60.68874, 62.27511, 63.83315, 63.99326, 64.79602, 67.61703,
    69.67011, 71.57149, 74.70484, 79.48899, 88.54491, 95.8951, 95.05336,
    95.01968, 95.02678, 93.84657, 89.89708, 82.89405, 79.62203, 72.85831,
    66.3242, 70.54633, 73.7272, 77.16171, 77.82213, 78.61967, 87.63425,
    82.10217, 56.51526,
  68.30836, 71.70788, 74.77542, 78.14034, 80.66331, 85.65406, 94.73337,
    98.13049, 97.49873, 96.93616, 96.59428, 91.818, 84.08336, 84.45701,
    84.96853, 85.45985, 84.95919, 80.21073, 75.03056, 73.54752, 70.06597,
    69.07957, 71.96957, 75.17227, 75.9599, 74.2422, 77.14978, 81.42281,
    70.02851, 50.48948,
  75.93668, 79.59022, 82.59845, 85.76808, 87.69278, 93.38971, 96.71603,
    84.3279, 76.0649, 74.80401, 71.32312, 67.7907, 65.89938, 66.58746,
    67.76992, 69.93197, 71.51528, 70.70787, 68.45364, 68.33663, 68.25053,
    69.44015, 72.06516, 74.02041, 73.39885, 74.43459, 79.10368, 76.6957,
    62.65172, 50.45178,
  76.43987, 77.73141, 78.59409, 79.17067, 80.42685, 80.88644, 71.91927,
    68.191, 69.20983, 69.36343, 69.25992, 69.53714, 71.62995, 76.49517,
    79.19753, 75.47672, 76.93135, 78.74871, 77.84011, 74.6028, 73.31386,
    76.64587, 80.30484, 79.7413, 77.74245, 82.75608, 83.367, 71.47329,
    52.86495, 51.221,
  81.60774, 84.33899, 80.94821, 81.84055, 83.96735, 80.00747, 67.09833,
    72.57258, 73.74009, 77.05975, 80.16753, 83.42979, 83.37926, 82.70778,
    81.45374, 84.22766, 85.51635, 84.58915, 82.73432, 81.57211, 81.91437,
    79.83961, 77.28922, 74.30887, 78.49982, 85.34753, 78.20142, 59.14593,
    50.60423, 50.35125,
  84.97537, 85.68884, 87.30775, 87.13692, 90.62638, 84.9301, 77.87902,
    81.79131, 84.99525, 85.31081, 78.6454, 69.72158, 69.00527, 69.68967,
    70.4519, 71.89444, 73.16754, 73.47277, 73.72089, 75.38004, 79.13554,
    76.34303, 69.82857, 68.99945, 74.03381, 73.38924, 60.20036, 50.95133,
    51.39399, 50.29634,
  98.15398, 93.0732, 100.0955, 103.0085, 95.99889, 83.88923, 84.23013,
    77.98833, 72.9236, 71.90825, 68.2651, 66.08157, 68.09477, 68.34283,
    66.74534, 67.41425, 67.06355, 67.45309, 67.82533, 69.91826, 74.22608,
    73.7478, 69.14226, 74.28313, 76.58693, 65.30045, 51.53691, 53.73502,
    51.98819, 50.87989,
  109.2955, 111.4426, 112.8338, 111.7842, 109.0942, 104.9361, 93.29327,
    80.87217, 87.02577, 79.29058, 75.50876, 73.69153, 78.15268, 80.30032,
    75.30579, 66.59195, 68.31106, 68.4704, 68.77989, 71.34613, 74.20889,
    73.68173, 71.28091, 67.89577, 65.47263, 59.77594, 53.22321, 54.404,
    53.36689, 51.77393,
  107.5921, 108.0622, 107.0394, 103.9225, 101.6885, 100.7987, 100.5238,
    99.98463, 97.94945, 97.72159, 97.39024, 95.84585, 95.85082, 95.65128,
    90.88441, 79.58656, 76.37699, 80.78787, 82.67184, 78.35812, 73.40878,
    69.26082, 64.65, 58.35535, 54.89265, 54.12072, 52.88336, 52.20058,
    52.09476, 51.41141,
  98.6664, 93.2974, 92.87751, 91.25809, 91.63814, 95.51752, 101.1641,
    99.42088, 94.37816, 93.94283, 91.16893, 87.41115, 87.57927, 89.60127,
    88.81586, 86.93616, 82.36686, 79.46249, 77.83002, 73.5063, 64.64349,
    61.8256, 56.72495, 54.05792, 54.11444, 53.69247, 52.54773, 51.61853,
    51.00073, 50.67271,
  84.03858, 85.72597, 86.28622, 85.28062, 84.12434, 85.26884, 86.73969,
    83.79366, 79.75137, 77.09091, 76.46445, 74.13186, 73.84148, 77.12752,
    75.3322, 74.36761, 73.96999, 69.71281, 67.05608, 62.9987, 57.55329,
    57.02668, 54.1808, 53.55006, 53.85968, 53.52115, 52.49321, 51.67405,
    50.98466, 50.62138,
  73.70415, 72.48846, 72.38718, 72.72253, 73.25754, 73.64629, 74.40682,
    75.4683, 74.59934, 72.42581, 69.81961, 72.97066, 77.33289, 75.03368,
    71.26807, 69.03091, 66.93491, 65.24471, 64.75601, 62.4634, 57.39532,
    57.36732, 54.68339, 53.62714, 53.56803, 53.44263, 52.21406, 51.09889,
    50.74326, 50.54563,
  66.6191, 67.22597, 66.9007, 68.0966, 68.86484, 70.16788, 71.3886, 72.87723,
    74.0296, 73.09863, 75.89046, 78.69157, 78.0895, 77.41783, 73.53728,
    70.11824, 66.35635, 65.93148, 66.66943, 63.28562, 57.23651, 56.65802,
    54.9401, 54.26271, 53.20688, 52.58693, 51.91428, 50.69817, 50.4911,
    50.36938,
  75.96965, 71.82294, 65.9305, 63.25911, 64.62243, 64.80519, 65.88605,
    67.3857, 67.88988, 69.43069, 72.3164, 71.74692, 68.45901, 69.78597,
    69.75078, 71.54334, 76.34863, 80.43167, 79.41159, 72.92513, 63.31745,
    57.99065, 55.40376, 54.6081, 53.15964, 52.28415, 51.67677, 50.76577,
    50.43479, 50.35836,
  75.47337, 70.62796, 64.76731, 61.30069, 62.41813, 62.93636, 64.09161,
    65.55332, 67.68932, 70.90823, 71.69958, 68.47569, 69.10799, 68.89143,
    68.18134, 68.9469, 71.88513, 75.27043, 75.28323, 72.65447, 66.90249,
    60.83324, 57.07886, 56.09012, 54.58247, 52.86311, 51.92365, 50.8869,
    50.42499, 50.38279,
  72.4198, 68.94544, 63.26209, 60.43792, 61.46329, 62.12652, 63.16579,
    64.55704, 66.60764, 68.67739, 67.20817, 64.604, 66.76, 66.47791,
    65.10933, 64.37919, 65.00826, 65.67528, 65.79491, 64.24868, 62.98898,
    62.01059, 59.90011, 58.02805, 55.74425, 53.45708, 51.84723, 50.91591,
    50.46778, 50.39748,
  70.98148, 67.92624, 62.4617, 60.12513, 61.03312, 60.58107, 61.39718,
    62.10951, 64.08109, 64.79796, 61.88185, 59.95841, 61.16259, 61.09431,
    60.74173, 60.89104, 61.23809, 61.73019, 62.01129, 62.07832, 61.97866,
    61.41253, 61.24622, 59.75122, 56.98215, 53.95406, 52.25059, 51.3347,
    50.6139, 50.39812,
  70.4221, 68.55213, 62.14099, 60.06378, 62.00642, 62.34536, 61.63183,
    60.20428, 60.61897, 60.01633, 57.59804, 57.92717, 58.84451, 59.4937,
    59.5323, 60.4343, 61.18768, 60.8188, 60.50019, 60.25434, 60.04379,
    59.61116, 58.86157, 58.35741, 58.28411, 55.85721, 53.29999, 52.45896,
    51.35831, 50.48995,
  73.99826, 73.27773, 68.93894, 67.39468, 67.67043, 66.54384, 66.59028,
    66.3531, 68.0684, 66.49217, 64.31993, 66.20441, 67.59531, 68.23745,
    67.49229, 67.12419, 66.78786, 65.24561, 62.95666, 61.47054, 60.5499,
    60.03328, 59.05222, 58.13425, 58.6301, 58.8627, 56.64663, 53.61622,
    52.48991, 51.09129,
  77.49502, 74.95735, 68.76514, 66.26064, 66.29052, 65.70198, 66.52089,
    69.09985, 72.53583, 70.26727, 67.53879, 70.02921, 72.02404, 72.43163,
    71.42998, 71.15134, 70.06127, 68.5205, 66.12029, 64.17212, 63.09875,
    61.87865, 59.97301, 58.53383, 59.11049, 60.45953, 59.92166, 56.14339,
    53.83966, 52.13153,
  80.0815, 78.52715, 72.44723, 67.82996, 67.0889, 66.98767, 69.69775,
    73.34866, 73.77296, 70.31031, 70.07619, 72.14912, 73.97419, 73.231,
    71.36593, 71.14324, 70.63802, 69.44337, 67.79643, 66.03216, 64.89615,
    63.2442, 60.57687, 59.20241, 59.64037, 59.90429, 60.22264, 57.25395,
    53.25802, 51.76075,
  80.39699, 77.91438, 72.64837, 69.02595, 68.1358, 67.1746, 70.07689,
    71.99872, 71.24053, 69.72997, 70.83936, 72.44441, 73.74438, 73.06042,
    71.87772, 71.5175, 70.99617, 70.06241, 68.84521, 67.96114, 67.86,
    67.75412, 66.04025, 64.00619, 63.41804, 63.16127, 63.29629, 60.09305,
    53.689, 50.86785,
  79.9319, 78.43027, 75.30032, 74.30121, 74.94559, 73.81568, 73.47953,
    72.46374, 70.21633, 70.56993, 71.77332, 73.72963, 75.40431, 75.89067,
    75.61755, 74.89664, 73.70354, 72.94299, 72.46004, 72.07726, 70.6795,
    68.04539, 65.48175, 64.28582, 64.05549, 64.05402, 63.53279, 62.73421,
    58.91524, 52.43674,
  71.08134, 71.29057, 72.28331, 73.23881, 75.17424, 76.58992, 73.31231,
    68.36954, 66.86008, 67.22937, 67.13593, 68.00967, 69.54335, 70.92922,
    71.72989, 71.45268, 70.33642, 69.00483, 66.69553, 64.37107, 62.99873,
    61.71112, 60.1477, 58.98497, 59.22412, 59.4672, 58.7894, 57.27223,
    56.17611, 53.31729,
  66.97667, 67.57767, 68.0965, 68.31314, 70.51553, 74.44439, 74.4683,
    68.2778, 65.53032, 67.00167, 67.77697, 68.60274, 68.8461, 67.98685,
    66.72842, 65.21515, 62.39179, 59.94043, 59.06276, 57.69491, 56.52455,
    56.33596, 56.30365, 55.99662, 55.82043, 56.02839, 55.31329, 53.82667,
    52.22686, 50.66587,
  46.91346, 46.89404, 46.90937, 46.89823, 46.89684, 46.986, 47.15593,
    47.44144, 47.70443, 47.98616, 48.57143, 48.4734, 47.39809, 47.58943,
    47.63646, 47.33166, 47.32533, 47.45266, 47.73148, 48.23602, 48.3633,
    47.84011, 48.16043, 49.4591, 50.8789, 51.10052, 52.03678, 53.1351,
    49.10774, 47.52268,
  47.80692, 47.82549, 47.62218, 47.83791, 47.70016, 47.73166, 48.04284,
    48.39666, 48.73616, 49.04495, 49.37378, 49.66812, 49.66444, 48.8404,
    48.28043, 48.40025, 47.98065, 48.2263, 48.77941, 49.25961, 49.24824,
    49.61468, 51.58529, 56.05575, 59.96062, 56.48864, 51.69373, 53.95349,
    49.64086, 48.02232,
  48.05196, 47.96585, 47.96181, 47.93397, 47.88018, 47.96245, 48.13846,
    48.42145, 48.63424, 48.8078, 49.0396, 49.29007, 49.55235, 49.91424,
    50.07467, 49.62482, 50.22466, 51.47737, 52.92008, 55.58028, 60.36206,
    66.51733, 69.40308, 68.46475, 66.6373, 61.52684, 57.83552, 53.36619,
    49.84766, 48.67795,
  48.69136, 48.86507, 49.46914, 50.0607, 50.45751, 51.07098, 51.33951,
    51.31031, 51.47921, 51.90331, 52.15162, 52.57249, 52.88743, 53.12487,
    55.0021, 56.76514, 57.17352, 58.09098, 61.94701, 67.25209, 74.16956,
    74.8036, 69.21886, 68.74932, 64.68208, 62.98186, 62.11635, 55.45093,
    49.424, 47.76497,
  51.2654, 51.46153, 52.39352, 53.05564, 53.19223, 53.22168, 53.2767,
    52.8717, 52.74611, 52.41321, 51.99685, 52.76578, 54.12069, 56.01553,
    58.43725, 61.36807, 62.8562, 63.64346, 67.48035, 72.50759, 71.82404,
    63.39498, 60.38391, 62.8335, 63.93055, 63.68837, 64.11511, 70.06287,
    68.28699, 54.42997,
  52.68979, 53.17703, 53.96131, 54.28793, 53.15998, 52.4915, 53.34267,
    54.28851, 56.17909, 59.59535, 64.85387, 74.66438, 83.6585, 83.5681,
    86.24303, 86.57438, 85.2894, 82.11638, 76.7769, 73.06781, 65.18163,
    57.5485, 61.39325, 64.60542, 68.17467, 69.59299, 71.57133, 81.48377,
    77.19128, 52.77127,
  53.74302, 55.11393, 57.07697, 59.35876, 61.53325, 66.75555, 77.12227,
    87.76578, 88.55035, 88.7101, 88.88448, 88.58598, 84.71452, 84.11971,
    83.41412, 82.47033, 80.8891, 75.15386, 69.43297, 66.77982, 62.93021,
    62.20935, 65.85212, 69.35379, 71.08366, 70.71627, 74.53109, 79.64628,
    67.01227, 46.83893,
  61.38869, 65.95463, 70.97221, 76.63458, 82.04004, 88.98667, 90.28041,
    89.91454, 85.45659, 84.21973, 79.71, 74.14458, 70.06786, 68.45993,
    67.28609, 67.49007, 67.41025, 65.45449, 63.2695, 63.33485, 63.57953,
    64.98318, 67.56845, 69.69142, 69.525, 70.79971, 75.5327, 73.47218,
    58.93321, 46.75382,
  74.4026, 79.23786, 82.45512, 85.3988, 89.08231, 89.60409, 81.22659,
    75.05555, 73.4288, 71.17955, 68.8279, 67.33921, 67.59549, 70.18442,
    71.23579, 67.65087, 68.15105, 69.33681, 68.9377, 67.25247, 66.85613,
    69.74258, 72.95229, 72.57912, 71.78583, 77.44589, 79.50704, 67.9101,
    49.43932, 47.36943,
  83.95544, 87.56644, 84.545, 85.0245, 86.44086, 80.54911, 66.17534,
    69.19633, 69.35811, 71.66568, 74.70683, 77.27554, 76.69659, 75.60094,
    73.97489, 75.34034, 76.18377, 75.4428, 74.2784, 73.98803, 74.74059,
    73.68104, 71.57928, 69.1103, 73.3105, 80.67118, 74.78165, 55.87355,
    46.92393, 46.87927,
  83.4086, 83.80676, 82.94505, 81.83054, 84.55731, 77.8485, 71.23305,
    76.3938, 80.57124, 82.3335, 77.11723, 69.27016, 67.71489, 67.41814,
    67.28336, 68.31171, 69.03388, 68.95749, 69.20555, 70.94452, 73.99911,
    71.86276, 66.8172, 66.54716, 71.91727, 71.33672, 57.65211, 47.32174,
    47.59958, 46.76693,
  84.90996, 79.11165, 85.77319, 91.41843, 88.36975, 80.87202, 83.7168,
    78.71591, 73.67759, 73.30229, 68.49026, 64.94224, 66.32564, 65.86363,
    63.78038, 64.3894, 63.77755, 63.83869, 64.04765, 65.57887, 69.26797,
    69.19978, 66.19028, 71.02463, 73.13914, 61.95285, 47.83036, 49.43877,
    48.19887, 47.17964,
  95.71791, 99.31217, 102.8565, 103.8041, 102.6045, 99.35925, 90.82606,
    77.39871, 82.29793, 75.50401, 71.16624, 70.1591, 74.08287, 75.26282,
    70.14072, 61.83586, 62.91535, 63.20865, 63.63921, 65.98604, 69.49698,
    70.54225, 68.95709, 65.19642, 61.75483, 55.4877, 49.17117, 50.55952,
    49.32162, 47.94173,
  101.8013, 104.5839, 104.2031, 100.7627, 97.45644, 94.66745, 92.76135,
    91.76391, 89.77085, 89.56993, 89.4658, 87.92003, 87.97273, 87.83726,
    84.07803, 72.33829, 70.364, 75.21599, 77.81883, 74.28658, 70.53284,
    66.52966, 61.39754, 55.26009, 51.26002, 50.30654, 49.31044, 48.75916,
    48.45749, 47.74514,
  99.36766, 98.12231, 95.42029, 92.62771, 91.06755, 91.86589, 94.10435,
    93.73237, 91.47244, 90.60487, 89.39258, 86.52145, 85.92637, 87.17789,
    85.95963, 84.38725, 80.29707, 77.95928, 75.89359, 70.44287, 61.25924,
    57.84369, 52.6909, 49.69626, 49.71743, 49.53224, 48.75164, 47.96486,
    47.44681, 47.07264,
  93.46898, 91.58554, 90.61938, 89.28291, 88.88889, 90.27109, 91.23451,
    87.76079, 83.34215, 79.47382, 78.01629, 75.78923, 75.63, 78.55624,
    76.43477, 74.42674, 73.06773, 67.72974, 63.74535, 58.91279, 53.69551,
    52.48621, 49.7635, 49.07483, 49.53569, 49.41353, 48.53424, 47.83379,
    47.27804, 46.98032,
  84.79895, 83.55621, 82.73614, 81.96587, 81.076, 79.3881, 78.65317,
    78.66306, 76.50385, 73.59317, 70.9716, 73.01125, 76.08338, 73.62969,
    68.8924, 65.93271, 63.12799, 60.43441, 58.83732, 56.54807, 52.57807,
    52.34997, 50.07508, 49.22743, 49.42208, 49.47475, 48.47956, 47.48424,
    47.12387, 46.974,
  76.21996, 76.04274, 74.76456, 74.51115, 74.00085, 74.05819, 74.29579,
    75.08816, 75.08685, 73.44644, 74.76086, 76.24036, 75.13015, 72.84328,
    67.71642, 63.91859, 59.99283, 58.81657, 58.9284, 56.50816, 52.44499,
    52.0904, 50.49224, 49.84758, 49.30301, 48.90389, 48.18872, 47.20018,
    46.96988, 46.83259,
  81.8178, 78.28107, 72.2924, 69.37318, 70.34529, 70.21773, 70.63382,
    70.94833, 70.10616, 70.06479, 71.10287, 69.02831, 64.77001, 63.68471,
    61.55534, 61.70978, 65.20892, 68.95772, 69.17931, 64.97029, 57.96537,
    53.5516, 51.15832, 50.48716, 49.42037, 48.6966, 48.08089, 47.17423,
    46.86245, 46.80266,
  81.33636, 76.3808, 69.74541, 65.85644, 66.36252, 65.94789, 65.88867,
    65.80546, 66.07837, 67.25386, 66.76514, 63.52415, 62.87773, 61.86179,
    61.01616, 62.10666, 65.54469, 69.27255, 69.3272, 66.55216, 61.52097,
    56.14668, 52.63667, 51.76107, 50.64701, 49.20604, 48.31706, 47.29063,
    46.81829, 46.81034,
  77.54467, 73.4913, 66.76839, 62.97968, 63.10565, 62.76159, 62.85756,
    63.33295, 64.5248, 65.76047, 64.47013, 62.89515, 64.75117, 64.61588,
    63.57098, 63.07857, 63.47707, 63.46424, 62.30279, 59.50384, 57.57928,
    56.5958, 54.82509, 53.18216, 51.51057, 49.69735, 48.27019, 47.36168,
    46.84338, 46.80214,
  75.35241, 72.08095, 65.73915, 62.68271, 63.13776, 62.74885, 63.47226,
    64.33125, 66.02905, 66.50411, 64.29347, 62.96295, 63.66875, 62.88248,
    61.4124, 60.21385, 59.10687, 58.30393, 57.44732, 56.62685, 56.26957,
    56.18985, 56.12186, 54.57818, 52.37222, 49.94858, 48.52331, 47.64308,
    46.96052, 46.82407,
  74.51982, 72.51369, 65.86073, 63.54657, 65.2692, 65.62119, 65.29166,
    64.47405, 64.79514, 63.48566, 60.61625, 59.96489, 59.6818, 58.94877,
    57.70062, 57.30408, 57.14563, 56.50317, 55.80966, 55.29239, 55.10344,
    54.94872, 54.31143, 53.39945, 52.94901, 50.92303, 49.11406, 48.4457,
    47.50115, 46.8912,
  76.06586, 75.4722, 70.59663, 68.88746, 69.24205, 68.07805, 67.49064,
    66.84663, 67.78913, 65.7762, 63.2425, 63.99243, 64.61492, 64.29543,
    62.85406, 62.02399, 61.5424, 60.1165, 58.00148, 56.52829, 55.51334,
    55.1132, 54.16196, 53.2875, 53.45686, 53.37703, 51.62349, 49.33481,
    48.41052, 47.33951,
  78.51274, 76.80563, 70.76491, 67.7105, 67.1591, 65.86699, 66.12083,
    68.07802, 70.96627, 68.63836, 65.8386, 67.53048, 68.53367, 68.19898,
    66.59322, 65.73701, 64.60625, 63.28947, 61.49408, 59.70617, 58.18102,
    56.78104, 55.06897, 53.93084, 54.47125, 55.31592, 54.63108, 51.37524,
    49.40364, 48.11365,
  79.59212, 78.30984, 72.22349, 67.39453, 66.31845, 65.66465, 67.66367,
    71.47304, 72.59119, 69.27223, 68.71517, 70.34383, 71.46739, 69.99036,
    67.6758, 66.73873, 65.91111, 64.83701, 63.39312, 61.6912, 59.93803,
    58.05658, 55.77227, 54.82383, 55.27914, 55.25439, 55.11279, 52.56286,
    49.26178, 47.865,
  79.74883, 77.89587, 72.71958, 68.74148, 67.74496, 66.67439, 69.02322,
    71.38936, 71.3287, 69.38985, 69.86604, 71.11042, 71.73438, 70.09234,
    67.83262, 66.77473, 65.63043, 64.30444, 63.03354, 61.99142, 61.59616,
    61.33675, 59.80784, 58.44292, 58.08108, 57.61278, 57.63303, 54.95885,
    49.53425, 47.21129,
  79.36692, 78.15861, 74.63562, 72.82703, 73.64724, 73.13789, 73.08871,
    72.62532, 70.42535, 69.76618, 70.13236, 71.24841, 72.20011, 71.50319,
    70.18251, 68.92622, 67.36684, 66.28127, 65.73589, 65.56342, 64.65604,
    62.66944, 60.41538, 59.22825, 58.99364, 58.59081, 57.94505, 57.2939,
    53.65826, 48.291,
  72.97038, 73.1974, 73.35306, 73.8763, 75.99413, 77.32591, 74.42534,
    69.88681, 68.03555, 67.79574, 67.17146, 67.34356, 68.25394, 68.82047,
    68.74621, 68.13621, 66.97786, 65.69815, 63.78004, 61.98487, 60.68394,
    59.1792, 57.55459, 56.43612, 56.30907, 55.77346, 54.72244, 53.37289,
    52.00098, 49.1586,
  68.67921, 69.19329, 69.50169, 69.6475, 71.64764, 75.02103, 74.82336,
    69.21572, 66.66566, 67.28886, 67.39844, 67.5947, 67.33802, 66.20906,
    64.71391, 63.04679, 60.50439, 58.1829, 57.06666, 55.66403, 54.45706,
    53.97259, 53.67554, 53.2386, 52.80937, 52.39237, 51.26376, 49.99195,
    48.78102, 47.25409,
  6.060241, 5.073979, 5.476762, 5.56749, 5.638362, 5.759594, 5.982664,
    6.274065, 6.725277, 7.613065, 9.348741, 11.5281, 13.36771, 17.02267,
    21.26226, 26.02434, 30.14175, 34.96923, 40.52453, 46.64471, 52.73629,
    57.75682, 61.46705, 63.88182, 64.99081, 64.95608, 63.24926, 65.40621,
    60.20452, 58.03192,
  4.578995, 3.819812, 4.123964, 4.621931, 4.883379, 5.106991, 5.476039,
    5.739035, 6.028511, 6.606508, 7.977128, 10.42784, 13.7661, 16.92615,
    20.91737, 25.19631, 29.99934, 35.40823, 41.28404, 47.84565, 53.77074,
    58.95316, 62.74095, 65.10601, 66.02079, 65.36298, 62.95653, 64.29309,
    60.36636, 58.59279,
  7.234473, 6.891779, 7.831794, 8.371229, 9.141071, 10.03453, 10.58853,
    10.67862, 10.84633, 11.25839, 12.11826, 13.59853, 15.90216, 18.93958,
    22.37149, 26.29762, 31.05606, 36.54982, 42.82061, 49.6152, 56.05912,
    61.36377, 65.04189, 66.71281, 66.89512, 66.28087, 65.79874, 64.93646,
    59.55998, 58.55698,
  9.852444, 9.869723, 10.29795, 10.28176, 10.41397, 10.53698, 10.65815,
    10.77788, 11.11473, 11.82692, 13.06931, 14.65729, 16.73629, 19.66741,
    23.27898, 27.22485, 31.83021, 36.80673, 42.97022, 49.82518, 56.52912,
    61.74517, 64.91682, 66.99775, 67.24, 67.16867, 67.11509, 66.17368,
    64.93418, 59.31845,
  11.37399, 10.36393, 10.85556, 10.82996, 10.89527, 10.8512, 10.89013,
    10.94736, 11.30616, 12.20191, 13.68537, 15.80188, 18.2641, 21.19595,
    24.6742, 28.62401, 33.1553, 38.28628, 44.27454, 51.17653, 57.14099,
    61.43348, 64.75232, 66.58521, 67.07189, 66.99682, 66.77249, 67.54018,
    67.19026, 65.27045,
  11.20434, 10.44299, 11.06272, 11.28846, 11.40224, 11.39684, 11.59814,
    11.76692, 11.82803, 12.28114, 13.53444, 15.64757, 18.68242, 21.84005,
    25.51545, 29.85703, 34.99697, 40.22702, 46.01065, 52.59166, 58.05818,
    62.03699, 65.24546, 66.58624, 66.79846, 66.4874, 65.97508, 66.55824,
    66.53986, 63.0638,
  11.1865, 10.35511, 10.98485, 11.22241, 11.52966, 11.8183, 12.23175,
    12.68125, 13.07482, 13.51557, 14.38755, 15.66973, 17.27682, 20.46519,
    24.36318, 28.86992, 33.92115, 39.89342, 45.7873, 52.6476, 58.3876,
    62.73099, 65.55969, 66.96558, 67.08028, 66.44337, 66.19966, 66.26221,
    65.59055, 56.61116,
  11.95995, 10.78201, 11.29935, 11.37256, 11.53589, 12.02181, 12.43795,
    11.50036, 11.0372, 12.36467, 13.65989, 15.55282, 17.97712, 21.02682,
    24.75872, 28.85724, 34.02108, 40.00331, 46.3539, 52.86369, 58.77546,
    63.1749, 65.93772, 67.10866, 66.96455, 66.70892, 66.85458, 66.42653,
    65.02739, 56.94345,
  14.82111, 12.88851, 12.72459, 12.37681, 12.14632, 12.05939, 11.21095,
    11.22848, 11.6645, 12.52497, 14.06559, 16.17873, 18.66231, 21.91996,
    25.7258, 29.15267, 34.0553, 40.64626, 47.48769, 53.82766, 59.49134,
    63.8868, 66.34215, 66.96194, 66.66867, 66.97441, 66.8663, 65.74371,
    57.28919, 57.51283,
  19.718, 17.52886, 16.19825, 15.07849, 14.53128, 13.53804, 11.7583,
    12.03604, 12.13365, 12.80855, 14.37581, 17.15205, 19.99022, 22.39875,
    25.39823, 29.71404, 34.68552, 40.54649, 47.04909, 53.97268, 60.23568,
    64.37066, 65.85847, 65.7892, 66.19172, 66.57915, 66.16265, 63.52615,
    56.77552, 56.54469,
  24.27385, 21.52692, 21.57757, 19.31953, 18.22882, 16.44304, 14.85749,
    13.89946, 13.77874, 14.67523, 15.65176, 17.66072, 19.7569, 22.70519,
    26.30506, 30.13872, 34.87399, 40.34768, 46.41998, 52.92952, 59.83614,
    64.10263, 65.48145, 65.72079, 66.17727, 65.87757, 64.6512, 57.11196,
    57.68235, 56.63475,
  24.56414, 22.08329, 24.76687, 25.05768, 23.94865, 20.52165, 17.49693,
    14.59343, 13.46156, 14.22937, 15.61661, 17.71524, 20.87618, 23.52064,
    26.58969, 31.10603, 35.31884, 40.84959, 46.9274, 53.02292, 59.0067,
    63.74258, 65.19292, 66.0285, 66.29981, 65.4133, 57.46003, 61.3055,
    58.14941, 57.27545,
  15.26194, 16.25561, 18.54263, 21.36419, 23.46543, 23.15029, 17.35598,
    12.31551, 15.81801, 14.8476, 16.55735, 18.01673, 20.55842, 23.42756,
    26.86876, 30.36782, 35.48007, 41.11741, 47.32913, 53.69674, 59.36261,
    63.2607, 65.03389, 64.99258, 64.99316, 64.69247, 58.05266, 59.54129,
    59.02919, 58.00401,
  11.83033, 10.45895, 10.60904, 10.84414, 11.44118, 12.2809, 13.29114,
    14.44884, 13.35683, 14.62804, 16.71067, 19.14212, 21.38601, 23.78045,
    27.33815, 30.98373, 34.888, 41.36707, 47.98748, 54.26555, 59.02594,
    62.53664, 64.10327, 60.66011, 57.76593, 58.00256, 57.55815, 57.17525,
    57.39258, 57.4651,
  12.62185, 11.39733, 11.98001, 12.01052, 12.3297, 12.50116, 12.84637,
    12.97609, 13.45286, 14.92498, 16.94283, 19.37263, 21.91271, 24.7541,
    27.33444, 30.68661, 35.60021, 39.80412, 46.87719, 53.64, 58.16866,
    61.8098, 60.64397, 58.8306, 59.27975, 58.49525, 57.745, 57.25734,
    56.79162, 56.73371,
  10.18808, 10.75101, 11.36324, 11.61435, 12.0829, 12.61575, 13.28681,
    13.65524, 14.31838, 16.22139, 18.93292, 21.21487, 23.56463, 25.46962,
    28.17691, 31.66326, 35.26827, 39.85535, 46.61542, 52.2854, 54.37372,
    58.74286, 59.05917, 58.98689, 59.08024, 58.57454, 57.75964, 57.25739,
    56.83326, 56.74147,
  7.36852, 5.729478, 7.345023, 8.862069, 10.67896, 11.40759, 11.97444,
    12.76304, 14.05636, 16.18349, 18.71503, 21.84707, 25.45518, 27.87209,
    30.65993, 33.6007, 36.94128, 41.73522, 48.36227, 53.80014, 54.79473,
    58.89587, 59.45321, 59.13241, 59.02061, 58.64685, 57.71152, 56.87112,
    56.61316, 56.66599,
  10.48071, 7.284759, 6.386683, 6.727334, 8.004313, 9.193612, 10.5327,
    11.55192, 12.46225, 13.96546, 16.79411, 20.34366, 23.75889, 28.54988,
    32.61718, 35.81641, 39.35021, 44.67656, 51.16722, 56.66137, 57.90622,
    59.40165, 59.72753, 59.69926, 59.00488, 58.39857, 57.71803, 56.76355,
    56.48835, 56.5406,
  22.33086, 16.09462, 9.259353, 4.302469, 6.257626, 6.44276, 7.432299,
    8.452571, 9.638637, 11.87822, 15.4176, 18.03114, 20.58229, 25.55813,
    31.10165, 35.76479, 40.99799, 47.62109, 54.9495, 60.58971, 63.42042,
    63.44185, 61.42392, 61.19616, 59.79572, 58.91727, 58.08887, 56.93853,
    56.46756, 56.58299,
  21.97657, 16.62853, 9.538216, 4.701846, 6.10809, 6.303149, 7.202435,
    8.330494, 10.22682, 13.29875, 15.68886, 16.16513, 19.34895, 22.20944,
    26.24307, 31.54661, 38.72645, 45.68735, 53.01099, 59.12156, 63.44693,
    65.54786, 63.42083, 62.58688, 61.04221, 59.40228, 58.39042, 57.12526,
    56.42907, 56.59803,
  22.75668, 18.09597, 11.44174, 6.733339, 7.684128, 7.581171, 8.262811,
    9.184047, 10.89865, 13.05604, 14.29599, 15.61605, 19.96113, 23.07437,
    26.44256, 31.06098, 37.10365, 44.41103, 51.76262, 57.95803, 62.62793,
    65.58752, 65.63895, 63.94571, 62.12216, 59.99904, 58.43353, 57.16161,
    56.4317, 56.59486,
  23.691, 19.59405, 15.12979, 11.19619, 12.70294, 12.16234, 12.73458,
    13.15896, 14.80346, 16.22532, 16.32939, 17.9449, 21.56461, 24.97099,
    28.45548, 33.04821, 38.56884, 44.93427, 51.36728, 56.75666, 61.14259,
    63.79923, 65.39111, 65.40145, 63.71466, 60.88823, 58.91872, 57.65843,
    56.6152, 56.5793,
  24.17786, 20.59276, 16.49755, 14.33284, 15.83792, 16.38256, 17.10858,
    17.75822, 18.86665, 20.18466, 21.86086, 24.59748, 27.69674, 31.07323,
    34.68489, 38.82086, 43.7872, 48.81007, 54.05412, 58.45181, 61.8872,
    63.94151, 64.75485, 65.15677, 65.53374, 63.15738, 60.12558, 58.56774,
    57.37503, 56.69857,
  24.17775, 20.36735, 16.8184, 15.13824, 16.45217, 17.04975, 18.31233,
    19.90706, 21.77247, 23.23103, 25.47655, 29.30253, 33.59572, 37.33906,
    40.44605, 44.35177, 48.8899, 53.92244, 58.91135, 63.54685, 66.16267,
    66.87814, 66.30119, 65.90587, 66.32123, 65.98838, 63.44452, 59.94197,
    58.45251, 57.41826,
  23.70367, 19.2967, 15.77481, 13.56508, 14.7765, 15.40187, 16.7395,
    18.73257, 20.7915, 22.26331, 24.5334, 28.58374, 33.28881, 37.33939,
    40.52923, 44.60908, 49.06926, 54.00991, 59.21381, 64.20337, 67.76733,
    69.164, 67.49261, 66.02782, 66.16927, 65.97494, 65.04839, 61.70402,
    59.1995, 58.26429,
  25.38189, 21.31692, 17.86353, 15.59423, 16.42181, 16.94865, 18.42368,
    20.41372, 22.1113, 23.55276, 26.20075, 29.98245, 34.4978, 38.21644,
    41.19098, 45.13266, 49.38631, 53.97385, 59.09521, 64.1517, 67.78603,
    69.54037, 69.35599, 67.93795, 67.66431, 66.62312, 65.79577, 62.91519,
    58.87366, 57.86413,
  34.55692, 30.88098, 27.52556, 25.21955, 26.11001, 26.39389, 27.7244,
    29.21087, 30.49975, 31.80407, 34.1492, 37.49702, 41.37609, 44.43921,
    46.72972, 49.84458, 53.02317, 56.56069, 60.70404, 64.99835, 68.22445,
    69.87155, 69.84495, 69.30634, 68.98016, 68.23805, 67.55494, 66.16673,
    60.57331, 57.36994,
  48.54864, 46.89548, 44.26178, 42.89392, 43.96702, 44.38303, 45.16165,
    45.8614, 44.75348, 45.6166, 46.97811, 49.45462, 52.15798, 54.13988,
    55.4402, 57.19295, 58.906, 60.62907, 63.20646, 66.07551, 67.88823,
    67.86551, 66.8882, 66.11823, 66.39272, 66.16763, 65.9249, 65.65063,
    63.55603, 58.78134,
  56.0181, 56.40978, 56.72431, 57.4804, 58.47184, 59.62981, 59.91526,
    58.05913, 56.59484, 57.02554, 56.73851, 56.81086, 57.27952, 58.0657,
    58.69495, 59.07589, 59.07492, 59.51526, 60.11012, 60.5493, 61.54684,
    62.66659, 62.72963, 62.10486, 62.27938, 62.25356, 61.62401, 60.10455,
    59.55642, 58.76579,
  60.63942, 61.32321, 61.59021, 61.67818, 63.03381, 65.11905, 65.7665,
    62.30258, 60.05203, 60.93568, 61.31623, 61.66862, 61.71902, 61.27753,
    60.81271, 60.30596, 59.18641, 58.05034, 58.10315, 58.21793, 58.05601,
    58.7736, 59.56895, 59.95097, 59.93028, 60.18544, 59.80533, 58.42774,
    57.49813, 56.80191,
  25.31098, 27.30712, 30.09304, 32.85149, 35.82361, 38.92281, 42.17515,
    45.56318, 49.10999, 52.65523, 56.20313, 59.45334, 61.97329, 63.93375,
    65.1697, 65.93636, 66.2773, 66.49203, 66.6601, 66.86305, 66.88367,
    66.69135, 66.54891, 66.51719, 66.28254, 65.51674, 59.90621, 62.70218,
    58.81581, 56.12349,
  24.24904, 26.20301, 29.17373, 32.33409, 35.35638, 38.86571, 42.60544,
    46.29199, 49.96414, 53.56665, 57.1035, 60.49951, 63.34956, 65.15097,
    66.0705, 66.53288, 66.67461, 66.8068, 67.01297, 67.33308, 67.64868,
    67.87166, 67.9632, 68.15211, 68.14065, 66.93015, 65.24709, 61.41969,
    58.11505, 56.48134,
  25.12433, 27.01269, 29.85518, 32.96535, 35.96933, 39.28699, 43.0527,
    46.95562, 50.86487, 54.54465, 57.91352, 61.05921, 63.78898, 65.74976,
    66.84582, 67.06867, 67.04061, 67.02152, 67.10731, 67.29485, 67.81281,
    68.39114, 68.58986, 68.60456, 68.37451, 68.04253, 67.38264, 65.69559,
    58.57681, 56.07346,
  25.85636, 28.01047, 31.26931, 34.122, 36.75026, 39.72002, 42.9827,
    46.97227, 51.06078, 55.13598, 58.7362, 61.76245, 64.41132, 66.28807,
    67.45985, 68.00934, 67.78441, 67.43062, 67.4753, 67.65308, 68.06574,
    68.07349, 67.48556, 67.86114, 67.65234, 68.0319, 68.39686, 67.74275,
    65.83409, 58.8037,
  26.52939, 28.88463, 32.00716, 35.37783, 38.17329, 40.84477, 43.61658,
    47.18278, 50.81866, 54.8455, 58.62564, 62.0609, 65.04429, 66.96848,
    68.24393, 68.90591, 68.80016, 68.19729, 67.88527, 68.03271, 67.88586,
    67.19939, 67.23421, 67.47933, 67.42165, 67.38803, 67.4996, 68.71096,
    68.34457, 65.70145,
  27.50591, 29.42873, 32.67053, 35.82096, 39.26052, 42.02546, 44.72478,
    48.31555, 51.53611, 54.66616, 58.18159, 61.75286, 65.07729, 67.07223,
    68.48551, 69.40685, 69.38332, 68.87984, 68.18859, 68.07529, 67.62801,
    66.88605, 67.44258, 67.62556, 67.5119, 67.28921, 66.92361, 67.57867,
    67.57198, 61.10613,
  30.71456, 31.42639, 33.70966, 36.39758, 39.479, 42.71467, 45.54595,
    49.25468, 52.77699, 55.71381, 58.68708, 61.29473, 62.89789, 65.16732,
    66.58687, 67.52724, 68.09315, 67.8776, 67.1564, 67.09164, 67.01548,
    67.05113, 67.39903, 67.72151, 67.7048, 67.42762, 67.28418, 67.28984,
    66.42741, 54.61221,
  35.71234, 35.61612, 36.71342, 38.3093, 40.56453, 43.68423, 46.81332,
    48.62297, 51.25502, 54.45756, 57.32483, 60.09751, 62.65944, 64.95386,
    66.5183, 67.36033, 68.07867, 68.39717, 68.02819, 67.449, 67.16353,
    67.16685, 67.41157, 67.62299, 67.40945, 67.5555, 67.69493, 66.97544,
    65.4503, 55.00141,
  41.45328, 41.96151, 42.09245, 42.52904, 43.5827, 45.48835, 46.65632,
    49.2586, 52.47065, 55.39822, 58.1525, 60.56868, 62.61653, 64.65959,
    66.47091, 67.04762, 67.66582, 68.5854, 69.1078, 68.60439, 68.00143,
    67.55445, 67.33617, 67.05326, 66.75163, 67.41451, 67.65578, 66.36172,
    54.8104, 55.49239,
  44.47721, 47.46216, 48.56857, 48.64023, 48.38868, 48.4527, 48.51561,
    50.77648, 53.41912, 56.46508, 58.93602, 61.24943, 62.97232, 64.21084,
    65.19936, 66.26199, 66.98361, 67.51611, 68.12855, 68.41286, 68.61266,
    67.84492, 66.97442, 66.25471, 66.46954, 66.7253, 66.45354, 62.07839,
    55.02319, 54.65503,
  42.97825, 46.32359, 50.96347, 53.30247, 53.92185, 52.8119, 52.46502,
    53.22272, 54.7319, 57.7783, 59.89578, 61.38852, 62.85415, 63.98894,
    64.91109, 65.64463, 66.23229, 66.58711, 66.95595, 67.25051, 67.97629,
    67.54578, 66.389, 66.40091, 67.0425, 66.52094, 64.51498, 55.79521,
    56.01532, 54.92752,
  39.16078, 39.64263, 47.17161, 53.13741, 58.3279, 57.56595, 55.21772,
    54.00105, 55.95015, 57.76773, 60.23043, 62.00512, 64.1532, 65.234,
    65.52184, 65.76942, 66.3699, 66.81347, 67.00655, 66.96948, 67.38312,
    67.23958, 65.92814, 65.94198, 66.65647, 65.99654, 54.9902, 59.95897,
    56.79659, 55.65977,
  33.28567, 36.06013, 39.42564, 45.54039, 52.39849, 57.49368, 56.00911,
    52.92121, 58.78356, 59.62176, 62.09246, 63.68294, 65.62207, 67.00263,
    67.18208, 65.91805, 66.46687, 67.17279, 67.50452, 67.18111, 67.2821,
    66.92475, 66.09204, 64.13809, 62.4844, 64.26434, 55.37921, 56.91806,
    57.1926, 56.29071,
  31.32312, 33.5946, 35.82476, 38.8336, 42.21188, 45.78223, 50.63615,
    55.68835, 57.16642, 60.23639, 63.17743, 65.59822, 67.09428, 68.21957,
    68.37556, 67.37811, 66.65677, 67.0955, 67.71455, 67.16664, 66.36388,
    65.92516, 65.16671, 59.86907, 55.40086, 55.43161, 55.61435, 54.89033,
    55.14339, 55.50502,
  29.53983, 31.09884, 34.64307, 38.46452, 42.09262, 45.72455, 48.94923,
    52.43661, 56.75522, 60.33847, 62.9851, 65.19528, 67.19344, 68.69826,
    69.02288, 69.16385, 68.21843, 66.97262, 66.54572, 66.24347, 64.4745,
    64.72673, 60.48018, 57.16116, 57.65638, 56.38404, 55.69533, 55.30299,
    54.85392, 54.78884,
  27.65503, 30.45697, 33.87335, 36.86359, 40.48952, 43.66715, 47.28848,
    50.84127, 54.73699, 59.03803, 62.39838, 64.95358, 67.16145, 69.08878,
    69.75792, 69.77622, 69.6486, 68.45972, 67.10925, 64.82954, 61.376,
    61.26633, 58.96321, 57.49756, 57.14076, 56.52626, 55.57069, 55.17568,
    54.96167, 54.88847,
  31.32685, 30.11557, 33.69481, 37.05721, 40.55594, 44.12271, 47.29148,
    50.12022, 53.46676, 57.22213, 60.67275, 64.07775, 67.14134, 68.78394,
    69.7607, 70.5899, 71.09644, 70.89277, 69.6702, 67.86044, 62.90625,
    61.82214, 59.78374, 58.08883, 57.38205, 56.71174, 55.67805, 54.88512,
    54.73395, 54.76564,
  39.48992, 37.00205, 36.27082, 38.17291, 42.46674, 45.46029, 48.83828,
    51.85853, 54.43128, 57.40265, 60.66948, 63.81757, 65.91117, 67.52807,
    68.50428, 69.62005, 71.01163, 72.11047, 72.3665, 71.01451, 68.34082,
    63.37601, 60.58813, 59.38958, 57.7963, 57.01392, 55.9689, 54.86328,
    54.66499, 54.70465,
  50.19717, 46.33693, 42.09643, 39.03114, 44.20969, 47.1892, 50.57999,
    53.93332, 57.12585, 59.88221, 62.64989, 64.80705, 66.19037, 66.84881,
    67.26317, 68.03644, 69.50792, 71.15208, 72.14592, 72.31953, 70.9985,
    68.27722, 62.4528, 61.24104, 59.10461, 58.05383, 56.74973, 55.17804,
    54.62144, 54.71209,
  50.05005, 47.65087, 43.47197, 41.82499, 45.76415, 48.63452, 52.39098,
    55.8541, 59.26167, 62.2273, 64.74476, 66.42439, 68.20583, 68.92153,
    68.92467, 68.121, 68.46398, 69.57613, 69.67817, 69.63213, 69.59234,
    68.79118, 64.99991, 62.7146, 60.64505, 58.76915, 57.16158, 55.43912,
    54.58728, 54.72918,
  51.4753, 48.78877, 45.18298, 43.83223, 47.83209, 50.71431, 54.47419,
    58.17989, 61.71635, 64.89135, 67.09997, 68.59168, 70.28333, 71.26841,
    71.41545, 71.29012, 71.13229, 70.99511, 70.51775, 69.13612, 68.5078,
    68.56847, 67.05303, 64.35783, 62.10248, 59.59849, 57.34277, 55.60815,
    54.63017, 54.73985,
  55.1193, 52.5598, 48.51431, 47.36115, 51.30263, 54.12441, 57.60174,
    61.08848, 64.79771, 68.29625, 70.85063, 72.55571, 73.80115, 74.32338,
    74.31528, 73.90292, 73.31245, 72.82395, 72.10881, 71.08585, 69.22655,
    67.48309, 67.02704, 65.7098, 63.92373, 60.69481, 58.13867, 56.45235,
    55.08767, 54.74878,
  62.04895, 59.19401, 55.06253, 53.35703, 56.7629, 59.286, 62.40285,
    65.45805, 68.6526, 71.84533, 74.83725, 77.50329, 79.1963, 79.58698,
    79.06832, 78.34358, 77.31649, 76.23721, 74.92131, 73.59695, 72.45545,
    69.88651, 67.56058, 65.97685, 65.73659, 63.11289, 59.51474, 57.56855,
    56.17742, 55.0083,
  70.74043, 67.2374, 62.77884, 60.7976, 63.11517, 64.52922, 66.91901,
    69.8215, 72.93988, 75.19346, 77.6902, 81.16127, 84.31441, 85.38483,
    84.26994, 83.65437, 82.41651, 80.68633, 78.55635, 77.23601, 76.09966,
    74.22837, 70.37142, 67.64906, 66.8904, 65.7647, 62.98603, 58.81038,
    57.12879, 55.98454,
  77.7156, 73.34908, 68.04327, 65.25214, 66.61718, 67.20046, 68.74866,
    71.15355, 73.89567, 75.3308, 76.86427, 79.67854, 83.12778, 84.51286,
    83.36306, 83.12919, 82.42788, 81.15925, 79.08717, 77.76577, 76.71297,
    75.01048, 71.79399, 68.72091, 67.76933, 66.38879, 64.79819, 60.70926,
    57.30776, 56.52974,
  80.76351, 76.1485, 70.84377, 67.67764, 68.23882, 68.18737, 69.5578,
    71.44615, 73.07458, 73.50771, 74.99965, 77.4598, 80.61961, 81.85536,
    81.00224, 80.86229, 80.46064, 79.45948, 78.2418, 77.32079, 76.10874,
    74.43957, 71.82391, 69.05979, 68.83549, 67.4081, 65.94733, 62.35261,
    57.52182, 56.06804,
  79.98133, 76.22919, 71.28511, 68.04665, 68.68388, 66.90913, 67.66601,
    68.97108, 69.3012, 68.73732, 70.298, 73.65481, 76.40841, 77.88763,
    77.37518, 77.59201, 77.29836, 76.57039, 75.61311, 75.12083, 74.38859,
    72.52624, 70.16096, 68.11168, 67.99742, 67.22803, 66.75378, 64.76638,
    59.34928, 55.92725,
  74.141, 72.19265, 69.15896, 67.2146, 68.16103, 68.1666, 66.73718, 65.84899,
    64.65569, 64.26784, 64.14636, 65.48678, 68.58079, 70.77278, 70.99317,
    70.92857, 69.82825, 68.69958, 68.22466, 69.01447, 68.93465, 67.82947,
    65.40752, 63.83951, 64.3506, 63.89286, 62.9509, 62.076, 60.57225, 56.99739,
  61.25879, 62.19572, 63.44622, 64.71423, 65.99062, 66.79277, 65.66003,
    62.0745, 60.8372, 61.1913, 60.61668, 60.07087, 59.9499, 60.7322, 61.106,
    60.93355, 60.14727, 59.54782, 59.09631, 58.80856, 59.3982, 60.52782,
    60.92374, 60.17668, 60.38789, 60.52261, 59.71879, 57.81482, 56.86843,
    56.46838,
  58.78905, 59.10379, 59.25027, 59.06023, 59.9174, 61.53554, 61.95472,
    59.4277, 57.83175, 58.57802, 58.86924, 58.87321, 58.63779, 58.24708,
    58.28846, 57.96895, 57.09012, 55.98199, 55.74579, 55.7005, 55.52637,
    56.17454, 57.07975, 57.55817, 57.4811, 57.71932, 57.55279, 56.38014,
    55.38339, 54.83797,
  60.85967, 62.60685, 63.63171, 64.67841, 65.29287, 65.76517, 66.0529,
    66.12139, 66.09157, 66.08775, 66.1083, 66.05833, 65.94267, 65.86013,
    65.71395, 65.59687, 65.5534, 65.41886, 65.31324, 65.08165, 64.54062,
    63.781, 63.18943, 62.77539, 62.40668, 59.69055, 54.61716, 56.91492,
    54.30577, 52.41837,
  60.73258, 62.55767, 63.57926, 64.70073, 65.39125, 65.9015, 66.23141,
    66.37965, 66.46925, 66.53454, 66.5095, 66.41875, 66.3527, 66.25266,
    66.03718, 65.88439, 65.70889, 65.5362, 65.49346, 65.47169, 65.2674,
    64.93983, 64.50833, 64.17288, 63.75359, 62.44325, 57.81276, 54.88287,
    53.82732, 52.64937,
  60.82696, 62.55043, 63.59922, 64.60033, 65.3082, 65.79332, 66.09524,
    66.33791, 66.56055, 66.72199, 66.74123, 66.63959, 66.47118, 66.43388,
    66.36506, 66.10806, 65.88583, 65.61864, 65.37335, 65.30654, 65.38668,
    65.3676, 65.13853, 64.88451, 64.29259, 63.50262, 62.69185, 61.02305,
    53.7182, 52.52906,
  61.02966, 62.74549, 63.72471, 64.66944, 65.36243, 65.91577, 66.2231,
    66.46341, 66.69108, 66.7556, 66.83993, 67.08169, 67.20109, 66.90096,
    66.73973, 66.65002, 66.32056, 65.89819, 65.74915, 65.51937, 65.47277,
    65.0198, 64.13672, 64.20104, 63.84918, 63.99141, 63.79852, 63.15934,
    62.1211, 54.7561,
  61.20802, 62.89462, 63.85326, 64.72401, 65.26176, 65.84261, 66.40437,
    66.62749, 66.64701, 66.5822, 66.6977, 67.40083, 68.0083, 67.77683,
    67.44653, 67.17948, 66.91318, 66.41547, 66.04025, 65.73151, 65.09012,
    64.26369, 63.72536, 63.65406, 63.62037, 63.49603, 63.52587, 64.36575,
    64.23644, 62.57204,
  61.75404, 63.1066, 64.15599, 64.8749, 65.31345, 65.86323, 66.58108,
    67.04224, 67.11783, 66.95207, 67.02789, 67.58058, 68.33223, 68.16572,
    67.96951, 67.70295, 67.11031, 66.70597, 66.22837, 65.7384, 65.02422,
    63.94828, 63.92773, 63.74087, 63.54472, 63.34087, 63.12595, 63.44915,
    63.57914, 57.94892,
  63.45506, 63.87378, 64.65971, 65.30457, 65.76856, 66.22926, 66.87212,
    67.07603, 67.15923, 67.19269, 67.28789, 67.00298, 66.29488, 66.49997,
    66.49043, 66.57629, 66.54078, 65.87505, 64.98971, 64.64966, 64.39394,
    64.0761, 63.98185, 63.97355, 63.81934, 63.61415, 63.52895, 63.43756,
    62.67893, 51.35188,
  67.24834, 66.28435, 66.19181, 66.37293, 66.65482, 67.17695, 67.36172,
    66.1551, 65.43004, 65.56481, 65.7181, 65.82188, 65.91914, 66.22493,
    66.54647, 66.68779, 66.73753, 66.42418, 65.6917, 64.95773, 64.3868,
    64.1597, 64.00994, 63.91371, 63.74959, 63.87433, 63.89588, 63.19662,
    61.96453, 51.58754,
  72.56089, 71.51595, 69.7952, 68.9187, 68.33261, 67.85739, 66.59412,
    66.47465, 66.3366, 66.06454, 65.86646, 65.64057, 65.49761, 65.71613,
    66.1781, 66.20852, 66.50826, 66.90065, 66.85355, 66.02384, 65.20625,
    64.45779, 63.97202, 63.417, 63.17685, 63.86795, 64.04428, 62.75217,
    51.51581, 52.10562,
  75.85318, 77.18198, 75.7512, 73.88351, 71.94157, 69.76067, 67.40298,
    67.34194, 67.16022, 66.94957, 66.19345, 65.64037, 65.15819, 65.00806,
    64.93688, 65.20344, 65.47101, 65.84803, 66.20483, 66.16997, 65.75645,
    64.84531, 63.91377, 63.04512, 62.9847, 63.17199, 63.04281, 57.86804,
    51.63475, 51.64404,
  74.26735, 76.96416, 79.76257, 79.24451, 77.37613, 73.42219, 70.53801,
    68.75795, 67.82207, 68.12845, 66.81793, 65.49554, 65.07728, 64.73869,
    64.45041, 64.44384, 64.48523, 64.00605, 64.44072, 65.08787, 65.32651,
    64.65342, 63.55738, 63.3512, 63.76266, 63.33858, 60.9819, 52.23132,
    52.69962, 51.73843,
  70.39455, 70.84536, 75.9929, 79.57845, 80.68764, 77.62846, 73.27743,
    69.86714, 68.7067, 68.31236, 67.60143, 66.66064, 66.40129, 66.07439,
    65.22987, 64.68906, 64.75958, 64.72936, 64.61785, 64.49838, 64.79322,
    64.43699, 63.26057, 62.92881, 63.23154, 62.90154, 51.98771, 56.69881,
    53.31384, 52.30086,
  64.62132, 66.62952, 68.3148, 71.59178, 74.94113, 76.38026, 72.06552,
    68.72504, 70.95121, 69.72135, 69.17812, 68.12508, 67.94823, 67.70253,
    66.77685, 64.9892, 65.06113, 65.22259, 65.0643, 64.49032, 64.52855,
    64.29133, 63.26208, 60.39221, 59.41481, 61.01259, 52.1897, 53.94588,
    53.8838, 52.9446,
  64.70248, 65.73414, 65.76154, 65.42674, 65.57339, 66.80762, 68.77705,
    70.15234, 68.84464, 69.74163, 69.9386, 69.19027, 68.68349, 68.37596,
    67.32871, 65.98975, 65.24993, 65.42474, 65.64931, 64.86761, 64.03875,
    63.34589, 59.54285, 54.99446, 51.76926, 52.05832, 52.37383, 51.747,
    52.03192, 52.33075,
  65.0382, 66.08495, 66.78011, 67.01646, 67.15643, 67.46124, 67.90932,
    68.03626, 68.16203, 68.16804, 68.27463, 68.17406, 68.41937, 68.29304,
    67.55402, 67.10535, 66.05688, 65.49362, 65.20084, 64.50005, 60.26538,
    59.92752, 56.20734, 52.91876, 53.69013, 52.97704, 52.41106, 52.10096,
    51.74614, 51.69912,
  65.24719, 66.66738, 67.23875, 67.49431, 67.43821, 67.77699, 68.04222,
    68.09889, 67.83472, 67.55417, 67.67804, 67.96354, 68.40571, 69.03728,
    68.48214, 67.66235, 67.28338, 66.38254, 62.90777, 59.99115, 57.57825,
    56.78625, 54.50408, 53.2984, 53.25062, 53.03334, 52.33555, 51.94893,
    51.80822, 51.76183,
  67.99944, 68.20825, 68.6596, 69.00708, 68.90508, 68.49824, 68.49276,
    68.66372, 68.35371, 67.90395, 67.60897, 67.99433, 68.91537, 69.21105,
    69.01626, 69.16057, 69.27545, 68.83833, 67.40152, 64.0376, 58.60748,
    57.44458, 55.31013, 53.87438, 53.66388, 53.25172, 52.29004, 51.69276,
    51.56688, 51.66072,
  74.08881, 72.20686, 70.6448, 70.41917, 70.71453, 70.44137, 70.2363,
    69.88419, 69.58176, 68.95273, 68.71734, 68.55514, 68.38759, 68.09325,
    67.85938, 68.6956, 69.87712, 70.49866, 69.99878, 68.22066, 63.59144,
    58.61148, 56.26752, 55.14406, 53.98011, 53.43464, 52.56283, 51.71344,
    51.54839, 51.57695,
  83.30645, 79.52259, 74.22556, 71.5099, 72.77466, 72.3332, 72.07024,
    71.49355, 70.8086, 70.43501, 70.35582, 69.95894, 68.0878, 66.06277,
    64.63087, 65.51212, 68.15865, 69.46889, 69.97256, 69.66464, 68.10877,
    62.87366, 58.04242, 56.99195, 55.20168, 54.29782, 53.2214, 51.95969,
    51.54068, 51.66964,
  82.93978, 79.91569, 74.75479, 72.46909, 73.90681, 73.93553, 73.82262,
    73.14883, 72.51459, 72.1673, 71.80387, 71.36365, 71.14106, 69.77827,
    66.54728, 64.80923, 64.57979, 65.828, 66.11198, 66.50369, 66.20425,
    63.91628, 60.07583, 58.2584, 56.45657, 55.03309, 53.66734, 52.1454,
    51.53874, 51.66789,
  82.4625, 79.56963, 74.8538, 72.36448, 74.04554, 74.52985, 75.06193,
    75.06049, 74.89496, 74.43555, 73.61974, 72.65594, 72.29593, 71.84689,
    70.94948, 69.63706, 68.48871, 68.00294, 66.73008, 64.24335, 62.96594,
    62.50621, 61.14546, 58.99385, 57.55418, 55.78343, 53.92791, 52.28705,
    51.51175, 51.65667,
  81.34035, 78.76628, 73.75054, 71.60239, 73.33771, 74.06631, 75.22031,
    75.94201, 76.77754, 77.24042, 76.55348, 75.21322, 74.37156, 73.83915,
    73.28594, 72.43365, 71.23512, 70.24521, 68.93679, 66.26158, 63.71815,
    61.69597, 61.59317, 59.72627, 58.62514, 56.71742, 54.78238, 52.99237,
    51.82186, 51.65019,
  80.06323, 77.64219, 72.66154, 70.55177, 72.409, 73.37858, 74.55141,
    75.7037, 77.43994, 78.8991, 79.1568, 78.66673, 78.31881, 78.06339,
    77.29829, 76.18265, 74.82388, 73.7632, 72.43472, 69.74268, 66.65159,
    63.9108, 62.36467, 60.56239, 60.34434, 58.54919, 55.843, 53.98979,
    52.6945, 51.81239,
  79.35194, 76.31216, 71.56844, 69.5372, 71.02837, 71.93269, 73.29335,
    75.157, 77.42022, 79.02067, 80.01959, 81.24821, 82.43533, 83.15376,
    82.11353, 80.92754, 79.41063, 77.52866, 75.88423, 74.0616, 71.76517,
    68.50641, 64.91426, 62.71007, 62.08455, 61.1007, 58.54575, 54.90434,
    53.54002, 52.63314,
  79.18301, 75.33236, 70.24841, 65.78712, 66.90028, 67.61105, 70.21908,
    72.95908, 75.62302, 76.57301, 77.55686, 79.0603, 81.51301, 82.30398,
    81.39636, 80.42952, 79.3186, 77.95, 76.22536, 74.84737, 72.97311,
    70.0955, 66.3148, 63.50418, 62.86186, 61.48609, 59.81741, 56.28097,
    53.66471, 52.9868,
  77.95721, 74.27094, 69.83978, 65.11092, 65.08385, 64.70609, 66.59277,
    69.83028, 72.3605, 72.58258, 74.08111, 76.01991, 78.5621, 79.75607,
    78.5722, 78.06734, 77.39145, 76.44216, 75.40559, 74.388, 72.70791,
    69.8884, 66.55409, 64.0641, 63.60148, 62.02839, 60.38823, 57.34944,
    53.77473, 52.5994,
  75.86125, 72.82225, 68.38114, 64.57854, 64.76576, 63.54476, 63.94254,
    65.11529, 66.01194, 65.70215, 67.58242, 70.79878, 73.84062, 74.82868,
    74.44005, 74.294, 73.68089, 72.93649, 72.39534, 71.84565, 70.33256,
    67.79398, 65.45151, 63.53284, 63.42976, 62.37951, 61.34321, 59.30397,
    55.21682, 52.72413,
  70.25665, 68.87916, 65.77312, 63.26166, 64.55946, 64.04922, 62.9251,
    62.18135, 61.2588, 60.82637, 61.01147, 62.3516, 64.9878, 67.25372,
    67.20609, 66.60815, 65.79654, 65.04471, 65.11885, 65.98849, 65.32834,
    63.82176, 61.46228, 60.23336, 60.43942, 59.8601, 58.88827, 57.83125,
    56.40326, 53.42339,
  57.26957, 58.46499, 59.48333, 59.92907, 61.08679, 62.77525, 61.2897,
    58.14791, 57.25695, 57.34311, 56.6326, 56.22453, 56.21619, 56.97934,
    57.11911, 57.05581, 56.32215, 56.04428, 55.68781, 55.74726, 56.28928,
    57.04372, 57.39197, 56.70929, 56.79736, 56.70684, 55.94924, 54.59703,
    53.72158, 53.0983,
  54.93087, 55.22197, 55.5864, 55.33532, 55.93111, 57.2917, 57.481, 55.65514,
    54.51427, 55.05365, 55.10725, 55.03973, 54.79374, 54.52151, 54.62697,
    54.30028, 53.6426, 52.76296, 52.62164, 52.52002, 52.42646, 53.02601,
    53.89966, 54.36141, 54.16976, 54.26383, 54.10997, 53.17968, 52.37187,
    51.83776,
  64.7087, 64.51067, 64.52105, 64.44921, 64.3155, 64.19659, 64.10608,
    64.05689, 64.03358, 63.77481, 63.51158, 63.56932, 63.40388, 64.08939,
    65.14213, 65.90373, 66.46846, 66.32988, 65.01012, 62.89494, 59.96221,
    56.41899, 53.73869, 52.09606, 49.98309, 46.49555, 43.92339, 45.53168,
    43.25084, 41.65156,
  64.57506, 64.42099, 64.42287, 64.40306, 64.19363, 64.02915, 63.99083,
    63.96357, 63.95088, 63.97509, 64.13197, 64.41994, 64.34213, 63.37759,
    63.04327, 63.71505, 65.23191, 67.4494, 68.42289, 69.45991, 70.41552,
    70.89977, 69.09547, 66.95497, 63.68968, 53.9201, 44.71354, 43.662,
    42.94639, 41.84461,
  64.62664, 64.58618, 64.67152, 64.61606, 64.4362, 64.25401, 64.18447,
    64.22353, 64.24463, 64.29543, 64.46381, 64.772, 65.14186, 65.5724,
    64.0649, 61.92204, 60.72036, 61.2261, 63.38766, 66.92506, 70.92606,
    71.95609, 72.24637, 72.13834, 69.93932, 65.02052, 60.19167, 46.60029,
    42.31343, 41.84341,
  64.53963, 64.5099, 64.71668, 64.74842, 64.62569, 64.48502, 64.43257,
    64.438, 64.47147, 64.4996, 64.73469, 65.22409, 65.69653, 66.01949,
    66.50649, 67.02699, 64.90859, 61.83471, 60.97585, 62.78483, 67.58864,
    67.29341, 59.92316, 62.81234, 62.57152, 69.17132, 70.70856, 64.34048,
    50.74276, 43.25461,
  64.50494, 64.41375, 64.6223, 64.6563, 64.58255, 64.64791, 64.88145,
    64.85119, 64.65466, 64.5713, 64.95919, 65.74795, 66.55879, 66.94984,
    67.3386, 67.90848, 68.17758, 68.18434, 68.70909, 65.48293, 61.74129,
    56.40969, 53.10645, 55.32295, 57.3175, 60.10085, 66.91948, 71.62251,
    71.73033, 52.63301,
  64.55623, 64.34903, 64.50854, 64.4108, 64.24152, 64.62359, 65.39713,
    65.67154, 65.42307, 65.07831, 65.19727, 66.06523, 67.09357, 67.4071,
    68.06719, 68.74313, 68.73868, 68.72586, 68.82126, 69.39413, 64.11318,
    53.08197, 56.18376, 55.39226, 55.32112, 55.02223, 55.65258, 63.99987,
    67.93062, 47.20332,
  64.96793, 64.49006, 64.46699, 64.27589, 64.16245, 64.59447, 65.47806,
    65.91626, 66.01337, 65.77441, 65.81573, 65.54873, 64.90054, 64.39485,
    62.66509, 61.52566, 63.02986, 61.7649, 59.01672, 59.09306, 56.93699,
    55.3398, 56.81955, 58.42763, 58.60867, 58.31229, 59.27096, 63.27135,
    58.25353, 40.78304,
  66.32623, 65.15939, 64.87773, 64.53474, 64.44553, 64.81665, 65.18887,
    64.25359, 62.63984, 63.89817, 64.1375, 64.01957, 64.24961, 64.41138,
    64.307, 63.52737, 62.26337, 60.48892, 58.33323, 56.40098, 55.46919,
    55.17394, 56.24773, 58.28255, 60.30849, 63.49389, 65.21337, 61.835,
    53.21147, 40.98261,
  69.59444, 67.69212, 66.4359, 65.63713, 65.1894, 64.8416, 63.82034,
    63.85926, 63.8678, 63.43458, 62.612, 62.3617, 62.56823, 64.23856,
    65.37847, 64.5106, 64.79447, 65.29606, 64.39413, 61.88789, 59.36787,
    57.73882, 56.88848, 56.37851, 58.31882, 65.63487, 70.77135, 60.04915,
    41.05027, 41.45794,
  73.77255, 72.53066, 70.61268, 68.77261, 67.52156, 65.93499, 64.09534,
    64.34177, 64.2848, 64.37402, 63.77926, 61.63096, 60.17581, 59.14419,
    58.6762, 59.53777, 60.57221, 61.78821, 62.71057, 63.09649, 63.06386,
    61.45752, 59.53516, 57.87457, 58.34667, 60.94572, 60.27981, 46.14878,
    40.95729, 41.03254,
  75.99647, 75.85648, 76.64172, 74.0602, 72.17917, 68.76579, 66.647,
    65.44281, 64.98901, 65.63294, 65.1335, 63.29676, 60.14487, 57.13308,
    54.98229, 54.53159, 53.82169, 53.78767, 54.59791, 56.40214, 59.09587,
    59.42688, 59.08743, 63.57789, 70.25523, 66.12264, 48.22735, 41.25844,
    41.74694, 41.10714,
  74.90536, 74.39792, 77.46483, 78.74991, 77.14702, 73.44248, 69.64794,
    66.44064, 65.07455, 65.48273, 65.32779, 65.0757, 65.57442, 65.80553,
    61.46378, 57.71022, 56.71286, 54.58973, 52.97344, 52.86243, 55.01219,
    55.67096, 54.36237, 56.7541, 63.00365, 60.26366, 41.52584, 45.16266,
    42.29113, 41.56298,
  67.11514, 68.70444, 70.54507, 72.96469, 74.94747, 74.73125, 69.28787,
    65.13128, 67.19837, 66.22746, 66.19342, 65.86044, 66.42252, 66.87829,
    66.73727, 61.7794, 63.0078, 62.4889, 59.64507, 55.84649, 56.28901,
    56.91986, 54.62779, 49.43001, 48.19247, 49.21275, 41.58281, 43.29768,
    42.98317, 42.11266,
  66.09639, 65.53329, 65.3269, 64.3927, 64.41455, 65.32298, 66.66525,
    67.28481, 65.78675, 66.29484, 66.67477, 66.58565, 66.65765, 66.96523,
    66.79893, 66.41128, 66.60414, 68.02328, 69.39348, 63.67244, 58.27534,
    54.05106, 46.8835, 43.77947, 41.24113, 41.49604, 41.63472, 41.23152,
    41.50499, 41.6236,
  67.55297, 67.27474, 66.76802, 66.0069, 65.53378, 65.66541, 66.22948,
    66.25352, 66.02431, 66.04411, 65.98241, 65.82056, 66.14416, 66.40491,
    66.27233, 66.37143, 66.48083, 63.17967, 59.0401, 54.27122, 48.1365,
    47.95218, 45.26261, 41.97054, 42.76342, 42.31258, 41.76085, 41.40403,
    41.17924, 41.15928,
  64.97895, 66.86542, 66.81759, 66.29905, 65.8514, 65.93034, 66.19826,
    66.44052, 66.37354, 66.37861, 66.56207, 66.62027, 66.8082, 67.10143,
    64.65855, 63.04079, 63.13821, 57.99788, 53.06721, 49.84793, 47.34842,
    45.56947, 43.14358, 42.22688, 42.38362, 42.37091, 41.7336, 41.33637,
    41.24163, 41.22111,
  66.09702, 65.24016, 65.22898, 65.40748, 65.29379, 65.13341, 65.76485,
    66.18818, 66.2043, 66.2868, 66.6379, 67.44387, 68.45724, 68.6211,
    68.11962, 67.04305, 64.1525, 61.14557, 56.62617, 52.47147, 47.97306,
    46.56779, 43.89676, 42.59916, 42.61751, 42.46084, 41.64828, 41.15251,
    41.10002, 41.14396,
  72.69485, 69.24477, 66.50565, 65.72253, 65.43902, 64.94314, 64.9698,
    65.20923, 65.34733, 64.85355, 66.04361, 66.93629, 67.74307, 68.30109,
    68.58089, 69.19033, 70.0554, 68.76942, 64.93758, 59.30573, 52.13332,
    47.62137, 45.04126, 43.69089, 42.96908, 42.54055, 41.77162, 41.129,
    41.10524, 41.1038,
  82.44363, 77.43937, 70.99075, 65.83061, 66.76922, 65.86649, 65.6745,
    65.22078, 64.07465, 63.53779, 63.33607, 62.08613, 59.60561, 58.50066,
    57.8853, 59.67091, 63.41319, 67.03621, 67.64276, 65.0541, 58.785,
    51.33859, 46.78689, 45.52913, 44.19381, 43.36822, 42.39182, 41.32463,
    41.06108, 41.15161,
  82.66909, 78.45802, 72.91897, 68.24292, 68.88758, 68.08269, 67.75612,
    67.15966, 66.72741, 66.64298, 65.8858, 64.21701, 62.92219, 59.01001,
    55.75846, 54.32726, 54.8838, 56.9528, 57.55676, 57.24725, 55.91025,
    52.46459, 48.31808, 46.61291, 45.18399, 43.95767, 42.76339, 41.45712,
    41.0463, 41.13177,
  82.4439, 79.37276, 74.04665, 70.65463, 71.57037, 71.02193, 70.79588,
    70.29324, 69.80624, 69.07377, 67.44384, 65.76579, 65.39858, 63.58788,
    60.84264, 58.99282, 57.6284, 56.72053, 55.23088, 52.78653, 51.49996,
    51.06581, 49.42495, 47.27402, 46.09814, 44.45514, 42.89767, 41.50532,
    41.02746, 41.16842,
  80.7401, 78.771, 73.58744, 71.62293, 72.86302, 72.96525, 73.20585,
    73.25141, 73.37347, 73.3484, 72.13508, 69.89034, 68.45622, 66.75877,
    64.70239, 62.88583, 60.87511, 59.14471, 56.83084, 53.50105, 50.72243,
    49.524, 50.45731, 47.92533, 47.27377, 45.31112, 43.58947, 42.03891,
    41.20041, 41.13453,
  78.98229, 77.52596, 72.48619, 70.606, 72.16396, 72.79556, 73.40302,
    74.09017, 75.40359, 76.42591, 76.51988, 76.16807, 75.7301, 74.51321,
    72.05265, 69.65073, 67.05482, 64.45602, 61.34848, 57.71545, 53.76025,
    51.2439, 51.02691, 49.01032, 48.97989, 47.19529, 44.82697, 43.08464,
    41.87162, 41.21913,
  77.0482, 75.0401, 70.95776, 69.21361, 70.4918, 71.18355, 72.18625,
    73.86362, 76.16224, 77.81496, 78.66264, 79.88667, 81.07891, 81.51566,
    80.35208, 78.88428, 75.46025, 71.43326, 67.86036, 64.0126, 60.3044,
    56.50182, 52.8542, 50.91636, 50.63483, 49.91814, 47.55871, 44.36354,
    42.82518, 41.89883,
  75.99853, 72.74711, 68.7179, 65.02331, 65.79848, 66.49075, 68.92429,
    72.22188, 75.08247, 76.29494, 77.21376, 78.79573, 80.80457, 81.47183,
    80.59696, 79.07671, 75.98246, 72.35033, 69.87302, 67.21782, 62.66447,
    58.38741, 54.02127, 51.35256, 50.94676, 50.16944, 48.6974, 45.5113,
    43.20906, 42.31281,
  75.39278, 72.15675, 67.77291, 63.22197, 62.98768, 62.85254, 65.08953,
    68.95461, 71.95738, 71.83282, 73.04974, 75.19189, 77.64142, 78.41248,
    76.85316, 75.36726, 73.20334, 70.92467, 69.31799, 67.24728, 63.30006,
    59.23711, 55.31177, 52.36433, 51.95171, 50.48694, 49.17536, 46.22035,
    43.139, 42.00938,
  74.72551, 70.15968, 64.20108, 60.48684, 60.19688, 59.08888, 59.94914,
    61.80435, 63.40487, 63.49507, 64.94423, 67.22176, 70.19434, 71.23122,
    70.36845, 69.34115, 67.41392, 65.74527, 64.87709, 63.85744, 61.16144,
    57.96988, 55.17083, 52.80978, 52.4393, 51.43384, 50.16847, 47.95734,
    44.20423, 42.00715,
  65.90715, 63.50731, 59.16902, 56.451, 57.26255, 56.39878, 55.56282,
    55.19499, 54.63699, 54.32382, 54.5735, 55.71211, 57.97651, 59.69025,
    59.43129, 59.05034, 58.2177, 57.34644, 57.09405, 57.326, 56.08476,
    53.86779, 51.26207, 49.92513, 49.96601, 49.34463, 48.32512, 46.95808,
    45.4537, 42.69644,
  49.71473, 50.46999, 50.99013, 51.24591, 52.16032, 53.54571, 51.66712,
    48.88187, 47.77022, 47.80307, 47.06293, 46.57709, 46.55988, 46.99585,
    46.93774, 47.09303, 46.82864, 46.66199, 46.49974, 46.53054, 46.74144,
    47.32957, 47.37362, 46.4239, 46.50554, 46.32083, 45.3956, 43.93199,
    43.13952, 42.44485,
  45.35214, 45.59606, 45.8079, 45.59571, 46.1937, 47.52185, 47.76469,
    45.60389, 44.44054, 44.88366, 44.95139, 44.86034, 44.52402, 44.21131,
    44.11765, 43.80413, 43.13886, 42.41846, 42.40296, 42.36484, 42.3175,
    42.96082, 43.82014, 44.14886, 43.878, 43.93021, 43.62934, 42.58938,
    41.86854, 41.32192,
  56.6634, 56.15931, 55.62232, 55.02997, 54.23622, 53.51313, 52.98818,
    52.71117, 52.76743, 53.2565, 54.18288, 54.98916, 55.14124, 55.82249,
    56.3571, 56.50623, 56.31846, 55.85374, 55.06416, 54.04487, 52.56348,
    50.70714, 49.84765, 49.98103, 49.45144, 46.4558, 44.36741, 45.7016,
    42.49083, 41.04768,
  59.97911, 59.57469, 58.85815, 58.29501, 57.32948, 56.37966, 55.55967,
    54.78291, 54.12975, 53.78123, 53.96956, 54.81379, 56.03187, 56.9434,
    58.10157, 59.78765, 61.27031, 63.02004, 63.46924, 62.3151, 61.30471,
    60.57018, 60.25684, 60.48095, 60.4904, 55.46267, 42.85385, 44.41782,
    42.35703, 41.3118,
  61.28416, 61.1698, 60.62372, 60.10502, 59.625, 59.32484, 59.06252,
    58.75645, 58.11668, 57.22207, 56.15359, 55.31739, 54.91057, 54.99398,
    55.38477, 55.77538, 57.43872, 60.30575, 63.84991, 63.01023, 62.44415,
    62.16718, 61.91146, 61.75195, 61.17405, 59.71027, 54.10964, 45.30513,
    41.82965, 41.47869,
  62.70798, 63.02391, 62.74308, 62.58817, 62.21884, 62.05853, 61.939,
    62.03056, 62.39814, 62.58163, 62.54499, 62.50148, 61.33407, 59.59206,
    58.88448, 58.09019, 56.89542, 57.28988, 60.48597, 63.39928, 62.75389,
    61.94831, 61.57574, 61.80595, 61.22462, 60.24934, 59.56096, 57.95894,
    47.18515, 42.2655,
  63.00929, 63.95295, 64.23753, 64.29664, 64.0765, 64.09711, 64.01249,
    63.00021, 63.01611, 63.72008, 65.77663, 69.85848, 70.29008, 69.59212,
    68.7715, 68.12114, 66.66459, 63.98252, 63.73345, 63.27939, 62.2098,
    56.10627, 56.47191, 60.60016, 61.00077, 60.57253, 60.40638, 60.91227,
    60.69368, 50.36218,
  61.77967, 63.48704, 64.55985, 65.52126, 65.78055, 67.61009, 70.79266,
    71.05532, 69.51865, 68.14195, 69.17018, 70.85532, 71.21793, 70.478,
    70.25804, 69.87086, 67.98341, 65.61745, 63.62715, 62.60484, 60.20001,
    52.19363, 55.96185, 57.41305, 60.39512, 60.77264, 61.00906, 61.64757,
    60.72048, 44.7653,
  60.97483, 61.94846, 63.17966, 64.54184, 66.00272, 69.93367, 71.39448,
    71.98193, 71.88391, 71.60931, 71.19543, 64.87376, 55.359, 56.04942,
    56.28368, 57.29556, 59.16555, 58.3701, 57.49507, 57.87881, 56.11568,
    54.8613, 56.65967, 58.45584, 59.47823, 60.52037, 61.08922, 61.19503,
    59.23084, 40.34721,
  63.54185, 62.73613, 63.33763, 64.24541, 65.99182, 70.29074, 71.20966,
    61.27075, 56.99413, 58.83778, 58.06367, 56.70129, 56.20665, 56.20272,
    56.22081, 56.2498, 56.3651, 55.91797, 54.81676, 54.45016, 55.0138,
    56.48201, 58.62457, 60.55804, 60.49842, 60.74651, 61.21329, 60.6637,
    51.2283, 40.50642,
  69.67043, 69.74818, 68.11923, 67.7698, 68.95285, 67.51488, 56.11272,
    54.6405, 55.46379, 55.50639, 56.40695, 57.2002, 58.0617, 60.59142,
    62.0136, 60.49063, 61.04119, 61.99483, 61.29248, 58.90704, 57.39315,
    58.16225, 60.03772, 60.45752, 60.50933, 61.14877, 60.85034, 59.27821,
    40.75183, 41.05159,
  72.92041, 72.8222, 72.31178, 71.92714, 71.47796, 69.89817, 55.8168,
    58.32307, 55.95691, 54.60055, 53.77977, 54.48685, 54.50293, 54.33652,
    55.00674, 57.25828, 59.21274, 60.54313, 61.32495, 62.09847, 62.6446,
    61.34783, 59.63054, 59.01639, 60.37781, 60.97077, 60.01842, 45.30244,
    40.47787, 40.48384,
  77.04279, 76.58058, 77.33575, 75.65216, 74.87398, 72.23935, 69.07268,
    67.17831, 65.25798, 62.51159, 55.47102, 50.31735, 49.38713, 48.79937,
    48.49506, 49.48722, 50.53099, 51.83809, 53.62876, 56.71933, 61.37368,
    62.00587, 60.3077, 59.92569, 60.25416, 59.81593, 47.43568, 40.63281,
    41.23661, 40.55374,
  81.30482, 80.20393, 82.40107, 82.67884, 80.21951, 76.77299, 73.49187,
    70.07928, 67.97462, 67.29044, 63.21985, 59.9205, 57.73426, 55.69395,
    53.05814, 50.61515, 50.64665, 50.30344, 50.2338, 51.65735, 55.80435,
    58.52913, 58.93093, 60.45849, 60.48508, 57.06504, 41.14498, 44.22308,
    41.76993, 41.04199,
  74.39412, 76.44128, 78.5293, 80.19481, 80.94403, 79.26777, 72.97734,
    69.26607, 70.21054, 68.37306, 67.48587, 66.69887, 66.40949, 66.54747,
    66.16877, 54.50106, 56.47846, 56.49675, 55.02607, 53.23104, 54.91458,
    56.58561, 54.8475, 50.71899, 50.27972, 48.15536, 41.40354, 42.98963,
    42.67087, 41.64004,
  66.53267, 64.95007, 63.95532, 62.71282, 63.84351, 69.46173, 71.02386,
    70.9566, 66.57287, 68.51525, 67.8836, 66.43768, 66.12394, 66.24123,
    65.36969, 63.54067, 61.90604, 63.62067, 63.35448, 62.1483, 57.97584,
    55.32701, 49.14929, 43.70625, 40.93886, 41.35756, 41.04963, 40.82282,
    41.13547, 41.10124,
  66.0088, 62.10426, 61.75605, 59.48121, 58.15979, 57.7714, 58.64755,
    58.25278, 56.55438, 56.39978, 56.4631, 56.3239, 58.90447, 59.67921,
    62.26281, 65.71268, 61.36351, 58.65352, 57.64297, 55.48042, 50.74451,
    48.13985, 43.65602, 41.74928, 42.30815, 41.85322, 41.26527, 40.89219,
    40.64786, 40.61161,
  59.175, 61.58106, 62.27192, 62.44794, 62.06467, 62.57788, 63.33732,
    62.15647, 59.41413, 56.81569, 56.16361, 55.29308, 55.11642, 56.63443,
    54.45743, 53.4377, 54.17817, 50.50589, 47.85267, 46.02025, 44.25723,
    43.99556, 42.20353, 41.65874, 41.97419, 41.93745, 41.27813, 40.9464,
    40.74987, 40.63643,
  56.05637, 55.80439, 56.25547, 56.9748, 57.67128, 58.30158, 59.56202,
    61.44785, 61.93044, 60.90852, 59.51211, 61.0376, 63.84387, 62.96822,
    57.90757, 56.12206, 53.68787, 51.84497, 49.57998, 47.51257, 44.43823,
    44.30128, 42.58855, 41.84089, 42.03265, 42.02486, 41.20727, 40.66989,
    40.63052, 40.62282,
  59.79246, 57.22742, 54.8929, 54.31254, 54.31928, 54.62466, 55.52717,
    57.09284, 58.56856, 59.33598, 61.40765, 63.39304, 64.66249, 65.57339,
    63.88321, 63.05442, 62.4499, 60.71117, 57.58458, 52.97919, 47.22689,
    44.91742, 43.38203, 42.59082, 42.10614, 41.77865, 41.18855, 40.59357,
    40.56329, 40.55622,
  73.74855, 66.72097, 57.86005, 52.83227, 53.28524, 52.3424, 52.31123,
    52.51424, 52.51655, 53.19008, 54.4268, 54.59089, 53.72712, 54.59404,
    55.36246, 57.55276, 61.79214, 65.29987, 64.99124, 61.60544, 54.7841,
    48.42103, 45.09115, 44.21264, 42.97962, 42.16139, 41.48833, 40.70848,
    40.50169, 40.56387,
  75.54126, 69.24832, 60.28157, 55.18404, 55.24935, 54.25563, 53.64583,
    53.12166, 52.96299, 53.39227, 53.04759, 51.52558, 51.4019, 49.79874,
    48.47052, 48.64263, 50.48932, 53.49616, 55.17561, 55.45179, 53.84755,
    50.36633, 46.88227, 45.3176, 43.98313, 42.7342, 41.77646, 40.8457,
    40.47794, 40.57249,
  77.91864, 72.75062, 63.8704, 59.02039, 58.92011, 57.76979, 57.05956,
    56.23947, 55.70821, 55.12266, 53.4496, 52.03323, 52.64259, 51.93996,
    50.48382, 49.91283, 50.10799, 50.91972, 51.29176, 50.46, 49.89811,
    49.70298, 48.16618, 46.50848, 44.96237, 43.29186, 41.99899, 40.93037,
    40.48484, 40.58887,
  78.42725, 75.54798, 67.35909, 63.34865, 63.67944, 62.50362, 62.07384,
    61.32865, 61.03903, 59.91564, 57.35814, 55.45507, 54.8299, 53.68242,
    52.34291, 51.7645, 51.39742, 51.5465, 51.54934, 50.96901, 50.34652,
    49.06187, 48.08504, 47.52334, 46.28128, 44.13481, 42.45304, 41.3404,
    40.60388, 40.57228,
  77.47983, 75.75284, 68.40698, 65.38646, 66.58766, 66.62396, 66.3422,
    65.86418, 66.41074, 65.81781, 64.15814, 63.60894, 62.69536, 60.90128,
    58.45997, 57.17873, 55.92897, 54.59196, 53.39172, 52.12284, 51.08076,
    49.57993, 48.12991, 47.98851, 48.08441, 46.04276, 43.5618, 42.19476,
    41.24488, 40.6645,
  75.15028, 72.72639, 67.40574, 64.99053, 65.58804, 65.40512, 66.12058,
    67.54315, 70.54617, 70.92413, 69.95296, 71.44261, 72.72542, 71.77689,
    68.83414, 66.84529, 64.46722, 61.69562, 58.9188, 56.51205, 54.5135,
    52.54611, 50.48329, 49.48944, 49.65734, 49.04122, 46.67376, 43.70156,
    42.34178, 41.26397,
  72.5938, 68.49393, 62.43201, 59.3918, 59.61445, 59.7267, 62.08013,
    66.02541, 70.04459, 68.97805, 67.79081, 69.1932, 70.82555, 70.89626,
    69.11058, 67.9262, 65.64825, 63.23428, 61.59228, 59.83478, 57.1688,
    54.6142, 51.80504, 49.77913, 49.7735, 49.21743, 48.13585, 45.07965,
    43.00943, 41.84456,
  70.21298, 66.66068, 61.18818, 57.11814, 56.48502, 56.33318, 59.32538,
    63.73499, 66.4342, 65.24716, 66.02182, 67.42266, 68.95132, 68.94092,
    67.40892, 66.37569, 64.73262, 62.93425, 62.09263, 61.05091, 59.08575,
    56.8781, 53.74763, 51.50528, 50.90659, 49.77834, 48.57208, 45.88357,
    42.72806, 41.5636,
  67.47148, 63.71694, 58.71746, 55.05136, 54.757, 53.75615, 55.56102,
    58.19883, 59.61879, 59.56163, 61.15295, 63.04287, 65.10108, 65.77369,
    64.87542, 63.8578, 62.15603, 60.70983, 60.27004, 59.78684, 58.63036,
    57.19765, 55.33838, 53.57758, 53.17009, 51.96268, 51.21507, 48.8592,
    44.11463, 41.33171,
  62.07268, 59.54341, 55.92805, 54.18902, 54.86707, 54.11176, 53.78016,
    53.58668, 52.75508, 52.97811, 53.80273, 55.33492, 57.3073, 58.21432,
    58.0606, 57.90599, 56.70567, 55.73762, 55.78638, 56.30384, 55.10632,
    53.29725, 51.21699, 50.1381, 50.46647, 49.99523, 49.33313, 48.76556,
    46.58266, 42.3996,
  49.31031, 49.96089, 50.44675, 50.94079, 52.4415, 53.95396, 51.93557,
    48.59634, 47.44677, 47.58575, 47.28163, 47.17213, 47.36432, 47.65623,
    47.46037, 47.57102, 47.32045, 47.04505, 46.73823, 46.75048, 46.91058,
    47.16011, 46.95174, 46.17249, 46.22882, 46.19176, 45.60394, 44.12986,
    43.45258, 42.40221,
  45.62681, 45.90476, 46.07432, 45.92865, 47.0603, 49.11011, 49.51772,
    46.2001, 44.74902, 45.53273, 45.80519, 45.96422, 45.80118, 45.2507,
    44.58966, 44.1607, 43.38247, 42.41017, 42.44711, 42.40442, 42.25491,
    42.82729, 43.60025, 43.85958, 43.69226, 43.82174, 43.48316, 42.27208,
    41.44819, 40.76967,
  50.95292, 51.23911, 51.57301, 52.01301, 52.36539, 52.87081, 53.40179,
    53.9802, 54.63838, 55.40087, 56.50717, 56.26114, 54.17553, 54.44971,
    54.8168, 54.72634, 54.89977, 55.49207, 56.08084, 56.88863, 56.67727,
    55.29721, 55.72676, 57.45794, 58.2076, 56.24827, 56.7286, 57.78138,
    49.36454, 46.64658,
  53.53151, 53.63641, 53.2764, 53.81517, 53.72317, 53.94037, 54.79883,
    55.7447, 56.8689, 58.12764, 59.71189, 61.33537, 61.56158, 61.43883,
    61.31838, 61.49449, 61.49006, 61.73517, 62.04215, 62.24396, 62.17071,
    61.99207, 62.00537, 62.56444, 62.75252, 61.43158, 53.38471, 55.98888,
    49.49356, 47.32335,
  55.7953, 56.07864, 56.15332, 56.13788, 56.0064, 55.97369, 56.08092,
    56.45535, 57.04773, 57.74046, 58.67577, 60.25658, 61.67723, 62.06786,
    62.28681, 62.11744, 62.15433, 62.46788, 62.81517, 63.23713, 63.70856,
    63.94491, 64.03575, 64.14294, 63.62936, 62.07352, 61.11384, 54.98763,
    48.95402, 47.82518,
  59.1846, 59.97842, 60.92688, 61.79904, 62.24752, 62.44532, 62.23104,
    61.97296, 61.83724, 61.63246, 61.55706, 61.92527, 62.13757, 62.03985,
    62.53242, 62.90721, 62.50508, 62.21241, 62.77838, 63.43818, 64.03673,
    64.09182, 64.35056, 64.97788, 64.39969, 63.00814, 61.7387, 60.95816,
    52.49921, 47.7033,
  61.9897, 62.78316, 63.66402, 63.29099, 62.79162, 62.48225, 62.43251,
    62.25511, 62.11759, 61.92765, 61.94727, 62.65012, 63.19435, 63.20318,
    63.33366, 63.86765, 63.49594, 62.40937, 62.55495, 63.24004, 63.27288,
    62.82588, 63.30502, 64.2178, 64.51937, 63.61346, 62.4103, 62.53277,
    62.40335, 56.08159,
  62.96423, 64.3656, 64.29734, 63.91496, 63.11401, 62.93433, 63.37285,
    63.15296, 62.66179, 62.37671, 62.61018, 63.55933, 64.46305, 64.34532,
    64.97215, 65.73238, 65.10374, 63.78973, 62.69033, 62.89145, 62.71113,
    62.33373, 62.91497, 63.51796, 63.9492, 63.72408, 63.13371, 63.67118,
    62.69983, 51.41961,
  61.97474, 64.53307, 64.52396, 64.25788, 63.54569, 63.61219, 64.35658,
    64.40754, 64.00365, 63.40822, 63.09936, 62.74851, 62.36857, 62.86594,
    63.5581, 64.19128, 64.16082, 63.19286, 62.30237, 62.68459, 62.75383,
    62.84714, 63.28926, 63.89606, 63.81693, 63.05064, 63.21266, 63.12621,
    61.48382, 45.78999,
  61.61775, 64.24148, 64.82626, 64.79555, 64.42829, 64.72991, 65.20261,
    64.31252, 63.57949, 63.55239, 63.38927, 63.37072, 63.50461, 63.80853,
    64.26558, 64.82439, 65.04443, 64.65401, 63.78305, 63.51083, 63.52892,
    63.96588, 64.59279, 64.77569, 63.97134, 63.57351, 63.86923, 63.15015,
    60.34079, 46.44523,
  65.77125, 65.62917, 65.36581, 64.95554, 64.29153, 64.18074, 63.95016,
    64.57776, 65.08516, 65.28168, 65.45089, 65.52736, 65.79898, 67.00378,
    67.68153, 66.62827, 66.94646, 67.42979, 66.98682, 65.57078, 64.7626,
    65.26975, 65.97588, 65.44003, 64.4429, 64.92173, 63.92533, 62.11562,
    48.02074, 46.83805,
  67.18334, 67.74381, 66.93053, 66.76947, 65.68295, 64.09949, 62.73597,
    63.53946, 63.88488, 64.66423, 65.14317, 65.49567, 65.2913, 65.03188,
    64.91194, 66.05818, 66.77844, 67.02901, 66.94954, 67.0064, 66.90971,
    65.48222, 64.03065, 62.68542, 63.36712, 64.18727, 62.65679, 54.08032,
    46.18557, 45.40139,
  66.87289, 66.7248, 67.87485, 66.58402, 67.17609, 65.34829, 64.22472,
    63.89901, 64.51782, 65.30864, 63.76495, 58.15413, 56.78526, 57.40004,
    58.11626, 60.21824, 62.67589, 63.08469, 63.59388, 64.70158, 66.42883,
    65.2151, 62.52883, 61.71544, 62.13707, 61.76799, 54.39751, 46.65586,
    47.06802, 45.55999,
  71.30631, 69.04079, 70.85196, 71.58896, 69.65825, 67.61125, 65.78243,
    63.39083, 61.85215, 62.48484, 62.21719, 61.32181, 62.12372, 62.64553,
    59.83268, 59.99711, 59.89989, 60.4451, 61.15653, 63.23278, 64.87189,
    64.82931, 62.59963, 62.82145, 62.59579, 61.07997, 46.98153, 50.79028,
    48.07397, 46.53457,
  70.76936, 72.08051, 73.46404, 74.5033, 74.05302, 71.94172, 66.09296,
    62.94101, 64.40854, 63.19047, 63.38405, 63.17471, 64.18748, 64.62685,
    63.09036, 62.08585, 62.28329, 62.60218, 62.84909, 63.55114, 64.26118,
    63.86862, 62.58291, 60.84594, 59.69937, 55.82751, 48.11016, 49.74393,
    49.55325, 47.6235,
  64.55206, 65.22366, 65.58474, 64.41047, 64.38067, 64.85, 65.69281, 65.8662,
    64.36538, 65.4872, 66.2144, 65.48933, 66.25351, 66.18504, 64.81684,
    63.1806, 62.54173, 63.18203, 63.75983, 63.65776, 63.33701, 62.67517,
    58.45906, 51.98909, 48.59287, 48.37953, 47.2674, 46.8463, 47.29247,
    46.88242,
  65.99722, 66.21517, 65.3393, 64.55585, 64.40562, 65.93292, 67.62407,
    66.00296, 64.42072, 64.23219, 63.89516, 63.27972, 63.68429, 64.45214,
    64.14334, 62.9848, 62.76469, 63.46981, 64.40136, 64.02888, 59.69207,
    57.22012, 51.71379, 49.72046, 49.92318, 48.84068, 47.59145, 46.75198,
    46.17348, 45.88213,
  66.11987, 66.51946, 66.29591, 65.52013, 64.89935, 65.27271, 65.75054,
    65.13082, 63.95384, 63.05059, 62.95481, 62.36054, 62.00089, 62.89644,
    62.53588, 62.10198, 62.64583, 63.08368, 62.69239, 59.17276, 53.29716,
    53.61022, 50.18773, 49.1919, 49.40654, 48.95602, 47.34481, 46.79221,
    46.31061, 45.88801,
  59.69666, 59.99454, 61.88324, 64.51253, 65.15187, 64.70702, 64.88928,
    65.62788, 65.39806, 64.66083, 63.67665, 64.24014, 65.40404, 64.43757,
    63.01848, 62.72464, 62.87955, 62.51047, 62.72401, 59.70236, 52.94707,
    53.92806, 50.9398, 49.27665, 49.06223, 48.83506, 47.03137, 45.93843,
    45.91165, 45.8065,
  57.40654, 57.15617, 56.87849, 58.76736, 60.78183, 63.19251, 64.693,
    65.32925, 65.82359, 65.59997, 66.1916, 66.94994, 66.92204, 66.85186,
    65.95146, 65.66097, 65.76718, 66.17012, 65.90009, 64.18043, 54.79816,
    53.60667, 51.51713, 50.2218, 48.3846, 47.55724, 46.91326, 45.69695,
    45.6745, 45.59601,
  67.72211, 62.12257, 55.34432, 52.28666, 54.45405, 55.46767, 57.50863,
    59.82907, 61.45993, 64.26286, 65.31258, 65.2737, 64.78153, 65.31665,
    65.47827, 66.6458, 69.01765, 70.88087, 70.41287, 68.37003, 64.82846,
    57.37514, 53.41895, 51.41383, 49.01217, 47.57705, 46.81367, 45.90963,
    45.61526, 45.60257,
  67.23651, 62.18687, 55.16252, 51.17709, 52.49358, 53.21902, 54.58649,
    56.22584, 58.60966, 62.29499, 62.8423, 58.93252, 59.93224, 59.73808,
    59.26052, 59.6722, 63.24528, 66.60435, 67.42098, 67.14792, 65.96018,
    61.75756, 55.95923, 52.7743, 50.61173, 48.36449, 47.0526, 46.05902,
    45.62243, 45.61425,
  68.04382, 63.51126, 56.24569, 52.25037, 52.62647, 52.86284, 53.80639,
    55.0956, 57.13411, 58.93926, 56.94381, 54.32897, 57.42642, 58.00173,
    57.37407, 56.84758, 58.00721, 60.0867, 62.43455, 63.0542, 63.26281,
    63.36944, 59.97258, 55.58807, 52.3541, 49.39613, 47.22265, 46.13215,
    45.59011, 45.61503,
  72.19135, 67.99699, 61.22008, 57.9423, 58.28833, 57.2805, 57.71405,
    58.07657, 60.11051, 60.34359, 56.31391, 54.65665, 56.34011, 56.68664,
    56.36648, 56.58406, 56.59166, 57.36566, 59.06409, 60.47879, 61.34243,
    60.64946, 60.30662, 59.37352, 55.80561, 50.74134, 47.8983, 46.85514,
    45.75589, 45.57094,
  76.15768, 74.6572, 67.46734, 65.18317, 67.15603, 67.34901, 66.33282,
    64.91733, 65.91134, 64.74596, 61.24855, 62.2232, 62.9252, 63.01816,
    61.93408, 61.48502, 60.77518, 58.90386, 58.44873, 58.93855, 59.22628,
    58.38496, 57.31635, 58.13174, 59.14058, 54.87775, 50.05545, 48.49307,
    46.93444, 45.71212,
  77.63522, 76.36279, 71.94306, 70.54608, 71.10951, 70.47079, 71.029,
    71.30107, 74.06499, 73.42211, 69.77986, 72.85773, 75.02219, 75.35661,
    74.19786, 72.55426, 70.59892, 67.59811, 64.24323, 62.70862, 61.78493,
    60.71359, 59.09327, 58.51492, 59.82135, 60.11901, 55.84812, 50.84611,
    48.80618, 46.71851,
  77.52833, 74.07548, 67.41353, 64.78545, 64.89695, 64.86805, 67.05532,
    71.41819, 75.51979, 74.08135, 70.1181, 72.93632, 74.86926, 75.91047,
    75.46149, 74.6379, 73.33414, 71.75047, 70.21613, 68.14633, 65.79828,
    63.30173, 60.46087, 58.54129, 59.03862, 60.09171, 59.47991, 54.19517,
    50.75797, 48.38543,
  78.23827, 75.70868, 70.97369, 65.75916, 64.09112, 63.67022, 67.72792,
    72.86262, 74.54273, 71.14621, 71.58626, 73.56382, 75.22417, 74.94757,
    73.77801, 73.72371, 73.42497, 72.71355, 72.35338, 71.65887, 70.61595,
    69.20592, 65.58345, 62.43972, 61.76811, 60.79045, 60.02005, 55.68056,
    49.48953, 47.57426,
  76.2767, 73.6527, 69.28491, 65.69931, 64.41087, 62.51614, 65.30912,
    67.9892, 67.68107, 66.74226, 69.04784, 71.21423, 72.86544, 73.20271,
    72.81438, 72.04078, 71.58633, 71.73498, 71.81374, 71.51794, 70.76205,
    70.13186, 68.88711, 67.76793, 67.18758, 66.30452, 65.4874, 63.01553,
    52.38497, 46.43562,
  71.32558, 69.7451, 67.32057, 66.24161, 66.87011, 66.62943, 65.93668,
    63.90141, 60.76988, 61.62564, 62.83525, 64.77361, 66.89468, 68.09519,
    68.84048, 68.30612, 66.91978, 66.70227, 67.87461, 68.81428, 67.06917,
    64.48456, 62.70779, 62.25198, 63.16988, 63.39317, 63.43792, 64.05595,
    60.01071, 49.36967,
  59.75475, 60.27098, 61.23159, 62.73474, 64.08745, 65.26968, 64.57901,
    59.27457, 56.99519, 57.99774, 57.45953, 57.60193, 58.41861, 59.54573,
    60.26722, 60.03479, 59.10442, 58.50117, 57.44396, 56.14597, 55.73158,
    55.49885, 54.51215, 53.69434, 54.45007, 55.00827, 54.56654, 52.83707,
    52.39493, 50.00065,
  55.07746, 55.51902, 55.62869, 55.64079, 58.65558, 63.93311, 64.56401,
    58.0937, 54.84799, 57.21037, 58.51746, 59.485, 59.38159, 58.964,
    57.76596, 56.35469, 53.08657, 50.35806, 50.08556, 49.65155, 48.78124,
    49.38871, 50.04386, 50.24801, 50.42222, 51.00423, 50.82026, 49.00574,
    47.13444, 45.70238,
  50.80473, 50.96244, 51.21502, 51.51244, 51.58468, 51.83491, 52.21806,
    52.70102, 53.35464, 54.40271, 56.69496, 56.59319, 52.71433, 53.2457,
    53.68726, 53.3121, 53.57932, 54.50085, 55.60213, 57.50343, 58.08078,
    56.45662, 57.27208, 59.92794, 61.87339, 61.60267, 64.94965, 65.23161,
    53.73196, 50.47211,
  53.88946, 54.33196, 53.64728, 54.50036, 53.98799, 53.68014, 54.22223,
    54.81801, 55.41027, 56.25766, 57.74793, 59.6909, 60.71063, 58.53967,
    57.11298, 57.92059, 56.99671, 58.27625, 60.1474, 61.69399, 61.38369,
    60.71061, 61.34411, 64.2923, 64.66421, 63.76324, 61.97297, 64.88277,
    54.89306, 51.62273,
  53.57507, 54.03893, 54.6735, 55.31607, 55.83459, 56.23431, 56.37985,
    56.78485, 57.33985, 57.97289, 58.84846, 60.33703, 61.92039, 63.97697,
    64.62157, 62.89425, 63.14654, 64.21271, 64.39865, 64.5007, 64.70958,
    64.89216, 65.02731, 65.53047, 65.55613, 64.40539, 64.23811, 64.48573,
    54.63877, 52.81352,
  56.26025, 57.08069, 58.56792, 59.90971, 61.23968, 62.91146, 62.89551,
    62.35079, 62.9276, 63.68144, 63.77989, 64.29738, 64.53114, 64.01452,
    65.09431, 65.62025, 64.8029, 64.10187, 64.52366, 64.94876, 65.39148,
    65.50711, 65.98357, 67.00616, 67.19041, 66.06682, 64.43164, 63.40292,
    55.79575, 51.21621,
  58.37794, 58.10511, 60.0961, 61.46256, 62.52955, 62.95097, 62.91204,
    63.08945, 63.79666, 63.80527, 63.84238, 64.62608, 65.18307, 65.37811,
    65.63705, 66.20787, 65.74278, 64.39879, 64.42176, 64.95324, 65.01792,
    64.66389, 65.25521, 66.57138, 67.6073, 66.4791, 64.05153, 63.92899,
    64.12857, 56.88357,
  60.75395, 62.82305, 63.58506, 64.08889, 63.77938, 63.65125, 64.31716,
    64.41074, 64.0005, 63.90198, 64.23288, 65.15757, 66.05299, 65.9865,
    66.61929, 67.676, 67.52768, 66.05679, 64.44284, 64.69714, 64.58136,
    63.86409, 64.96151, 66.0637, 67.04839, 66.37935, 64.58748, 65.1077,
    64.74295, 55.60612,
  62.57293, 62.98401, 63.69568, 64.12448, 63.90312, 63.98539, 64.51122,
    64.63479, 64.20811, 64.12685, 64.23144, 64.3429, 64.4103, 65.07745,
    65.80991, 66.59415, 67.17554, 66.15417, 64.49769, 64.90011, 64.88778,
    65.11803, 65.78495, 66.93375, 66.88863, 65.3304, 65.0117, 65.01712,
    64.2648, 50.84846,
  62.56969, 62.93127, 63.7014, 64.2467, 63.99224, 64.3256, 65.08878,
    64.52994, 63.81542, 64.02564, 64.20551, 64.55975, 64.88599, 65.58794,
    66.45914, 67.42506, 68.22303, 67.99265, 66.54913, 66.1201, 65.96593,
    66.46174, 67.51831, 68.08479, 66.87177, 65.87653, 66.33247, 65.9771,
    64.6298, 51.2547,
  64.33398, 64.55324, 65.12068, 65.08381, 64.34415, 64.79193, 65.35312,
    66.14809, 66.95266, 67.53381, 67.91785, 68.20982, 69.12588, 72.10871,
    73.85122, 71.39105, 72.05683, 72.99271, 72.3632, 70.27239, 68.80682,
    70.02238, 71.74651, 70.70257, 68.07174, 68.68714, 67.46771, 65.56979,
    55.1613, 50.92951,
  69.20029, 70.6512, 70.33806, 70.80239, 69.10294, 67.49297, 66.41016,
    67.5829, 68.43748, 70.28259, 71.86636, 73.25717, 72.94802, 71.64854,
    70.35416, 72.25904, 73.57355, 74.09265, 74.17841, 74.50043, 73.80413,
    72.06188, 70.1287, 67.58849, 67.14876, 67.16444, 65.84557, 59.48295,
    50.73549, 48.46574,
  67.67242, 67.35705, 68.8185, 68.58815, 69.58043, 69.17864, 68.61273,
    68.73219, 69.85591, 70.37918, 68.61682, 64.9509, 64.65894, 64.76854,
    65.04381, 65.58231, 66.46262, 67.1259, 68.19671, 69.34551, 70.883,
    69.92547, 65.50504, 63.72699, 63.94525, 63.80472, 56.91402, 50.93811,
    50.44318, 48.60224,
  71.16885, 68.65897, 71.62877, 72.26335, 70.8849, 69.68109, 68.67858,
    66.69433, 64.75289, 64.40855, 63.99629, 62.77943, 63.88495, 64.72551,
    64.69267, 64.46315, 64.43861, 64.86779, 65.34377, 66.66618, 69.26294,
    68.71711, 64.71901, 64.96107, 64.55745, 62.67843, 51.29994, 53.24503,
    51.6927, 49.74178,
  74.91112, 76.4563, 78.26996, 78.20956, 76.93109, 73.84441, 67.34534,
    64.82597, 66.06587, 64.05067, 64.43752, 64.11372, 65.06216, 66.05768,
    65.82925, 65.09684, 65.43939, 65.89908, 67.14819, 69.10944, 68.70338,
    67.42861, 65.0139, 64.36807, 64.12847, 59.10587, 52.61776, 53.38322,
    53.39064, 50.82517,
  68.05466, 68.72705, 69.17982, 68.07848, 67.51633, 68.07622, 69.29304,
    69.42575, 66.85211, 66.92476, 67.36849, 65.84446, 67.12174, 67.90382,
    66.60363, 65.64509, 65.56271, 65.87532, 66.62981, 67.1502, 66.44759,
    65.28712, 64.41766, 58.44568, 55.07998, 54.0997, 51.72089, 50.7907,
    51.23794, 50.36267,
  64.64074, 65.37021, 65.93803, 66.06631, 65.99051, 66.93849, 69.70893,
    70.1813, 67.83478, 67.51469, 66.87407, 66.57767, 67.33472, 67.51381,
    66.75684, 66.31997, 65.96933, 66.67253, 68.09618, 68.03066, 63.57503,
    62.44455, 57.67657, 56.40144, 55.75948, 53.65646, 51.89995, 50.75017,
    49.86063, 49.18571,
  65.30647, 66.08346, 66.87734, 66.84006, 66.77655, 67.98553, 69.61428,
    69.14361, 67.87323, 66.95931, 67.2286, 66.21531, 65.35919, 66.80125,
    66.34261, 65.96095, 66.55241, 66.85719, 67.61951, 66.77757, 58.17375,
    59.00953, 55.43875, 54.86272, 55.19027, 54.37058, 51.75655, 50.79332,
    49.93126, 49.15134,
  64.18166, 63.85282, 64.423, 65.00778, 65.59016, 65.79894, 66.80739,
    68.10449, 68.09593, 67.47008, 66.15876, 67.42861, 69.84599, 68.25577,
    66.41167, 66.14864, 66.29298, 66.59441, 67.53582, 66.88328, 57.50361,
    59.44907, 56.22964, 54.43895, 53.59093, 53.32553, 51.17072, 49.4299,
    49.33751, 49.04464,
  63.84877, 64.14806, 64.2432, 64.90038, 65.37478, 65.96218, 66.43243,
    66.80972, 66.95534, 66.60538, 68.07021, 70.32726, 70.08617, 68.77853,
    68.85954, 67.67647, 66.82906, 67.43001, 68.75396, 66.77418, 58.59614,
    57.82645, 55.95813, 55.00652, 52.55204, 51.62103, 50.90502, 48.89291,
    48.87119, 48.65273,
  68.42384, 66.61633, 63.86058, 62.12891, 63.6041, 63.67474, 64.1989,
    64.9243, 65.22532, 65.8485, 67.25969, 67.2485, 65.92697, 66.72322,
    66.87013, 67.95498, 70.31046, 72.52294, 73.38248, 71.36168, 66.90707,
    60.29438, 56.57655, 54.8238, 51.89678, 50.37783, 49.97965, 49.11037,
    48.7307, 48.62971,
  68.94102, 67.25171, 63.25285, 60.90067, 62.03483, 62.91268, 63.87472,
    64.66984, 65.44305, 67.09867, 67.71725, 66.0638, 66.17212, 65.97811,
    65.84962, 66.36922, 68.30525, 70.13931, 69.99841, 70.23182, 68.29693,
    66.10579, 59.24213, 56.41495, 54.07668, 51.2077, 50.1309, 49.19088,
    48.71646, 48.60954,
  66.14692, 64.7832, 61.48057, 59.24689, 59.4699, 60.18184, 61.14132,
    62.5315, 64.9389, 66.17957, 65.78108, 63.05742, 65.66525, 65.60138,
    65.00746, 63.16676, 63.88192, 66.10362, 67.25936, 66.74357, 66.73482,
    66.96252, 65.86311, 60.73599, 56.33667, 52.46482, 50.27052, 49.30396,
    48.73925, 48.63034,
  66.80953, 63.09097, 60.37383, 58.98456, 59.42946, 58.60247, 59.94665,
    61.31306, 64.90933, 65.61263, 61.82653, 57.89869, 60.94456, 61.888,
    61.5227, 61.93829, 62.28921, 63.00904, 64.89977, 66.00635, 66.06619,
    66.21806, 66.426, 66.1208, 60.88101, 54.08932, 50.88044, 50.01005,
    48.96972, 48.64296,
  67.10394, 66.07595, 62.29044, 61.70531, 64.85981, 65.22778, 65.03393,
    63.72604, 65.32287, 64.6534, 58.21225, 58.91195, 60.73279, 62.44154,
    62.21054, 63.35234, 63.98558, 61.95478, 61.47743, 61.43123, 60.86282,
    60.63754, 60.91737, 63.03648, 64.93166, 59.46994, 53.32211, 51.92055,
    50.52293, 48.83,
  70.2961, 69.17016, 66.63458, 66.13091, 66.46938, 66.43209, 66.98566,
    67.86201, 69.41818, 68.77473, 62.16845, 64.52345, 66.67901, 68.95248,
    68.67643, 68.6264, 69.05936, 67.31514, 63.98655, 62.41138, 61.10381,
    60.30154, 59.86842, 60.06982, 62.66501, 65.22266, 60.47984, 53.94981,
    52.31602, 49.68351,
  71.78501, 70.0574, 66.60436, 65.2002, 65.92316, 66.14104, 66.81353,
    68.65711, 71.29632, 71.08514, 65.05209, 66.78314, 67.73668, 69.00109,
    69.46893, 71.12212, 71.39188, 71.13039, 69.31936, 66.17724, 64.24815,
    63.29704, 62.25664, 61.25882, 61.71513, 65.03403, 66.44135, 59.94072,
    55.79456, 52.18338,
  72.7626, 71.19559, 68.4659, 66.32198, 66.17648, 66.24583, 67.93478,
    70.42989, 71.40012, 70.63875, 69.82656, 69.69476, 70.16406, 69.26514,
    68.52617, 70.24916, 71.18254, 71.2236, 70.88654, 69.97589, 68.75213,
    67.50369, 64.94011, 62.54757, 62.9733, 64.1059, 66.28496, 62.02285,
    54.42787, 51.53363,
  72.81699, 70.88314, 68.43472, 66.34624, 66.38528, 66.07597, 67.71748,
    69.35674, 69.48042, 66.957, 69.77244, 70.41429, 70.36754, 70.56747,
    70.91165, 71.32079, 71.70704, 71.8885, 71.76152, 71.22256, 70.44454,
    70.30672, 69.81582, 68.88206, 68.65884, 68.71674, 68.71116, 67.10979,
    57.32723, 49.3106,
  70.2821, 69.91893, 68.51039, 67.95052, 68.92156, 68.93768, 69.15095,
    69.1381, 66.61559, 68.48319, 69.5574, 69.64813, 70.14783, 70.67063,
    71.09133, 71.4241, 71.54302, 71.72161, 72.04519, 72.12706, 70.99057,
    69.87407, 68.98059, 68.49252, 68.57885, 68.46642, 68.26929, 68.20215,
    66.57693, 53.49738,
  65.54518, 65.4667, 65.87547, 66.37755, 67.94992, 69.351, 69.03449,
    67.05212, 66.07413, 66.70552, 66.58807, 66.90142, 67.37949, 67.63583,
    67.82509, 68.03611, 67.99107, 67.86938, 67.18118, 63.80513, 61.4388,
    60.37897, 57.9487, 56.71733, 58.39334, 60.4839, 61.20953, 59.77254,
    59.47226, 55.08594,
  65.00868, 65.30398, 65.50255, 64.87785, 66.54187, 68.96709, 69.80054,
    67.59481, 66.42787, 67.19328, 67.83904, 68.56635, 68.46954, 67.46145,
    66.44439, 66.00748, 63.4866, 58.60435, 57.5222, 55.93013, 53.84813,
    54.00262, 53.94858, 53.86433, 54.43386, 55.82854, 56.28147, 54.02073,
    51.07982, 48.68652,
  47.38342, 47.71051, 48.02396, 48.3663, 48.66193, 49.00891, 49.39317,
    49.87505, 50.43254, 51.12885, 52.8248, 52.79498, 50.5105, 50.91383,
    51.16843, 50.76261, 50.85096, 51.37739, 52.03855, 53.43048, 54.04076,
    53.22657, 53.85051, 55.33673, 56.00629, 55.31726, 58.22218, 58.30655,
    49.64203, 47.01039,
  52.51353, 53.15427, 53.16522, 54.18027, 54.29388, 54.60763, 55.3623,
    56.1139, 56.91049, 57.76672, 58.81417, 60.09975, 60.84503, 59.47624,
    58.66954, 58.84778, 57.901, 58.43848, 59.52309, 60.3499, 60.12352,
    59.56427, 59.92134, 62.57629, 66.20866, 63.98337, 60.36113, 61.16133,
    51.17778, 48.07702,
  55.18326, 56.08632, 56.96298, 57.97923, 58.92476, 59.90157, 60.88963,
    62.05273, 63.29219, 64.4155, 65.49915, 65.93389, 66.25786, 66.74551,
    67.28915, 67.65405, 68.27489, 68.89954, 69.19707, 69.22246, 69.28593,
    69.23431, 69.17307, 69.37402, 69.37239, 68.66286, 66.19732, 60.58162,
    51.67661, 49.31628,
  60.63718, 62.41968, 64.27019, 65.20416, 65.4585, 65.82658, 66.07037,
    66.17245, 66.31635, 66.31362, 66.33761, 66.88851, 67.22035, 67.14052,
    68.06105, 69.05962, 69.19856, 69.29603, 69.79741, 69.96004, 70.13254,
    70.1316, 69.98789, 70.79715, 71.08786, 69.70061, 68.33576, 59.22707,
    51.54609, 47.90135,
  65.32171, 65.46064, 65.79749, 66.08477, 66.08686, 66.40063, 66.9334,
    67.11388, 67.2035, 67.10783, 67.05455, 67.54958, 67.99435, 68.20394,
    68.58308, 69.42365, 69.64953, 69.47269, 69.85514, 70.25294, 70.45232,
    70.01223, 70.06727, 70.41303, 70.90649, 69.87303, 67.76279, 67.4392,
    62.91346, 51.225,
  66.17329, 66.58428, 67.06686, 67.28872, 66.8778, 66.96678, 67.72094,
    67.84055, 67.54937, 67.43691, 67.52803, 68.25101, 68.90869, 68.72528,
    68.98901, 70.3167, 71.76773, 71.18134, 70.10863, 70.2072, 69.8646,
    69.53385, 69.54339, 69.79541, 70.17315, 69.30978, 67.67585, 68.19189,
    68.24666, 49.97453,
  67.01072, 67.43465, 67.7777, 67.85055, 67.4328, 67.49685, 68.08493,
    68.17371, 67.70309, 67.5221, 67.51693, 67.49811, 67.41524, 67.54955,
    67.96423, 69.3894, 70.85586, 70.53141, 69.73276, 69.74867, 69.51346,
    68.45281, 69.11446, 69.99227, 69.82913, 68.34505, 68.12616, 68.37633,
    65.67957, 47.32936,
  67.25816, 67.54613, 67.75332, 67.85499, 67.38529, 67.27465, 67.745,
    67.37946, 66.73222, 66.73013, 66.79197, 66.83402, 66.94154, 67.27146,
    67.93536, 69.24405, 70.65848, 70.94911, 70.07306, 69.8204, 68.7793,
    68.80004, 69.93121, 70.20117, 69.40557, 68.75929, 69.19909, 68.86999,
    57.6735, 47.57977,
  68.53683, 68.78387, 69.03533, 68.93732, 68.42772, 68.57355, 68.82564,
    69.30846, 69.94094, 70.16235, 70.32851, 70.51604, 70.82635, 72.40641,
    73.47881, 72.60817, 73.52808, 74.42535, 74.11255, 72.78193, 71.8839,
    72.42534, 73.30302, 72.33733, 70.37439, 70.34621, 69.81796, 65.25764,
    51.16378, 47.29653,
  74.1345, 74.95947, 75.30087, 75.8632, 74.9189, 73.27789, 72.64357,
    73.48904, 74.06059, 74.80563, 75.22762, 75.95425, 75.85427, 74.93661,
    74.29056, 75.32543, 75.84153, 75.41177, 74.14983, 73.52074, 73.45476,
    72.66462, 71.49511, 69.76057, 69.7159, 70.6843, 69.27112, 52.12823,
    47.3574, 45.80076,
  76.80071, 77.59503, 79.21278, 79.31986, 80.54488, 79.25703, 77.86533,
    77.2098, 76.8624, 77.24818, 76.6945, 71.86602, 71.31115, 71.20734,
    71.67004, 72.39724, 72.94124, 72.62254, 71.9725, 71.54777, 72.09202,
    71.10526, 62.93481, 58.41382, 59.49444, 58.61612, 51.83094, 47.05544,
    46.58165, 45.74468,
  77.9482, 74.73226, 77.39289, 78.90844, 78.65813, 77.53287, 76.61226,
    73.87482, 71.00665, 70.55714, 69.70482, 68.41824, 68.62899, 69.25032,
    69.35101, 69.67656, 70.03448, 70.1329, 68.7291, 67.67592, 68.87157,
    64.5221, 56.93802, 61.37901, 63.23006, 52.11656, 46.96866, 47.5947,
    47.05482, 46.1736,
  82.32207, 82.60727, 84.12711, 84.88734, 84.0006, 81.02689, 74.19272,
    70.73896, 71.27448, 69.06108, 69.55611, 68.966, 69.21323, 69.57622,
    69.26988, 69.22538, 69.99162, 70.18054, 69.58192, 70.25868, 68.90334,
    61.61002, 57.52867, 57.96343, 57.96767, 50.63434, 47.83631, 48.01916,
    48.01482, 46.77802,
  77.97155, 78.42794, 78.422, 76.5103, 74.97514, 74.01987, 73.7858, 74.26989,
    71.99012, 71.83, 72.5611, 71.09151, 72.26111, 72.85926, 71.26945,
    70.44735, 70.57571, 71.08101, 71.14511, 70.67973, 67.95195, 61.36974,
    60.91542, 53.46179, 49.85883, 48.99166, 47.64915, 47.03521, 47.19475,
    46.57379,
  71.12687, 70.99828, 70.63447, 70.11, 69.99442, 71.17918, 74.74557,
    75.91055, 73.61564, 73.45995, 73.0261, 72.47205, 72.41212, 71.91548,
    71.09024, 70.26433, 70.52298, 71.05162, 71.79281, 70.87017, 62.02974,
    58.73579, 52.84698, 50.15881, 49.11514, 48.62474, 47.51927, 46.80062,
    46.47005, 46.08152,
  71.63966, 72.15283, 72.6031, 72.58092, 72.6068, 73.60648, 74.59403,
    74.5873, 74.20203, 73.30861, 72.7788, 71.20859, 70.15439, 70.62744,
    69.77418, 69.69053, 70.42151, 70.78343, 69.62981, 64.98725, 54.59332,
    53.51885, 50.90641, 49.84656, 49.25372, 48.58077, 47.53281, 46.8946,
    46.4869, 46.0267,
  71.74343, 71.79008, 71.91199, 72.08082, 72.64539, 72.56689, 73.04508,
    73.7593, 73.3508, 72.60502, 71.29148, 71.35703, 72.16559, 70.53124,
    69.40481, 69.50952, 70.29615, 68.73141, 69.25536, 66.39963, 53.66992,
    53.67517, 51.39908, 49.91568, 48.82825, 48.48018, 47.39525, 46.41433,
    46.23936, 45.99895,
  70.05396, 70.60967, 70.53401, 70.85085, 70.94466, 71.30054, 71.54454,
    71.94691, 72.3163, 71.46242, 71.54269, 71.87654, 71.09115, 70.37059,
    70.19762, 69.63813, 69.50944, 64.96848, 67.37662, 63.59218, 54.17913,
    53.0708, 51.07263, 49.59648, 47.87352, 47.50682, 47.00933, 46.10649,
    45.98352, 45.82756,
  71.97208, 71.11871, 69.77515, 69.03654, 69.47892, 69.43142, 69.84136,
    70.40851, 70.25326, 70.15438, 70.5882, 70.00758, 68.82089, 69.4222,
    69.94992, 71.14727, 73.11393, 74.25513, 74.56839, 72.85114, 61.27538,
    54.38715, 50.96994, 49.43404, 47.43854, 46.82513, 46.57884, 46.11294,
    45.92255, 45.80542,
  71.63558, 70.52798, 69.21168, 68.35734, 68.86161, 69.21377, 69.60609,
    69.91081, 70.19067, 70.89508, 70.85051, 69.56298, 69.6329, 69.91093,
    70.44313, 71.45695, 73.14699, 74.31913, 74.07826, 72.82638, 65.46882,
    57.55863, 51.89663, 49.86413, 48.12994, 47.03727, 46.56621, 46.18279,
    45.90554, 45.8026,
  71.03643, 70.2144, 68.81758, 68.10587, 68.52612, 68.91253, 69.32036,
    69.61895, 69.96323, 70.38762, 69.7294, 68.6841, 69.00134, 69.21501,
    69.53684, 69.72941, 67.66426, 66.59216, 66.6369, 65.35672, 63.21802,
    60.88395, 55.80686, 51.76114, 49.2513, 47.70702, 46.65065, 46.20958,
    45.93758, 45.81165,
  71.6021, 69.93529, 68.64127, 67.84533, 68.16616, 68.20914, 68.47606,
    68.60475, 69.01517, 68.97159, 67.81987, 67.14056, 67.24873, 67.40132,
    65.86022, 63.84203, 61.90861, 60.68537, 60.06456, 59.0627, 59.5774,
    60.11094, 58.74392, 57.49807, 53.07359, 48.93004, 46.9814, 46.56908,
    46.01885, 45.82261,
  71.21962, 69.85558, 68.29565, 67.42747, 67.84819, 67.90278, 67.55962,
    67.12879, 67.39603, 67.04747, 65.14051, 65.06497, 65.30924, 64.77449,
    63.12556, 62.07212, 60.69231, 58.21643, 56.9201, 56.35105, 57.04475,
    57.6953, 55.95499, 56.20976, 55.79713, 51.50768, 48.00963, 47.57003,
    46.65143, 45.89172,
  72.38584, 71.08097, 70.00466, 69.34932, 69.31111, 69.02559, 69.02216,
    69.29978, 69.73463, 68.82387, 67.44411, 68.22621, 68.68269, 69.209,
    67.36206, 65.16888, 63.375, 60.73666, 57.98115, 57.02744, 57.26075,
    56.87476, 55.32243, 54.28823, 54.53542, 54.33002, 51.02743, 48.35603,
    47.35178, 46.23199,
  73.79182, 74.14124, 71.70995, 70.71762, 70.84329, 70.72807, 70.64022,
    71.22845, 72.39481, 71.87742, 70.52281, 70.93273, 71.43508, 71.31961,
    68.82317, 66.66791, 63.97503, 61.78265, 59.17332, 56.74146, 56.45874,
    55.93032, 54.48027, 53.26342, 52.33054, 53.40213, 53.41954, 50.59667,
    48.8912, 47.23432,
  76.23524, 76.94566, 74.94386, 73.48223, 72.99703, 72.61922, 73.14889,
    74.08623, 74.03094, 72.92906, 72.11537, 72.19462, 72.52876, 70.92078,
    67.16605, 65.05183, 63.25398, 61.68063, 59.60375, 57.25856, 57.06343,
    56.71087, 54.5808, 52.88966, 52.47413, 52.71737, 53.68739, 51.97494,
    48.6487, 46.9983,
  77.19205, 77.60696, 75.48365, 74.10406, 73.86534, 73.39098, 73.74542,
    74.05512, 73.48509, 72.67999, 72.25, 72.17684, 72.23944, 70.36469,
    67.76535, 65.56876, 63.92222, 63.13133, 61.75465, 60.46277, 61.9641,
    64.03143, 63.11822, 59.44306, 57.02733, 56.20107, 56.79417, 55.2982,
    49.12913, 45.97946,
  77.22449, 77.28747, 75.70048, 75.07675, 75.4162, 75.01163, 74.45409,
    73.92245, 73.09344, 72.8783, 72.7077, 72.74613, 72.94563, 73.04951,
    72.62031, 70.59901, 68.56384, 67.87698, 67.45206, 67.36073, 67.81911,
    66.57197, 63.02472, 59.99873, 58.12169, 57.41246, 56.48872, 57.71731,
    54.69887, 47.61984,
  73.33176, 73.491, 74.47661, 75.12664, 75.52626, 75.79819, 74.87321,
    73.05621, 72.32024, 72.25639, 71.82759, 71.43681, 71.3318, 71.76264,
    72.61142, 73.31651, 73.45785, 71.56873, 67.74004, 63.76285, 62.01432,
    60.00391, 57.46508, 55.62522, 55.15073, 54.89166, 53.96715, 52.3452,
    51.79052, 48.83639,
  71.84871, 72.17085, 72.78532, 72.96596, 73.64864, 74.72598, 74.57743,
    72.67413, 71.53677, 71.69227, 71.59894, 71.30618, 70.95191, 70.7085,
    70.8116, 71.08845, 67.14416, 62.16116, 59.44057, 56.72186, 54.69341,
    53.81543, 52.98029, 52.19617, 51.6289, 51.49874, 50.88494, 49.29059,
    47.57726, 46.08158,
  38.58859, 38.69198, 38.78718, 38.87996, 38.90214, 38.9637, 39.06022,
    39.20586, 39.40901, 39.66787, 40.76208, 40.9062, 39.34673, 39.48468,
    39.65335, 39.26113, 39.18446, 39.44082, 39.72573, 40.60444, 41.09459,
    40.50833, 40.79392, 41.8368, 42.52637, 42.26415, 44.86991, 46.12971,
    40.93345, 39.21903,
  40.57209, 40.81197, 40.56326, 40.9557, 40.84229, 40.77008, 40.98479,
    41.19893, 41.42958, 41.70514, 42.14114, 42.76934, 43.20005, 42.21041,
    41.48744, 41.63163, 41.03907, 41.47341, 42.36061, 43.1847, 43.35476,
    43.29594, 43.89872, 45.4701, 50.30656, 51.1337, 45.54682, 47.80065,
    41.76519, 39.81465,
  42.65388, 42.90501, 43.02804, 43.24479, 43.41246, 43.60019, 43.76094,
    43.98954, 44.26882, 44.51302, 44.79803, 45.33638, 45.62671, 46.01662,
    46.00897, 44.84721, 44.85439, 45.72177, 46.36975, 47.35375, 49.13617,
    51.30774, 52.42306, 51.8259, 55.55087, 57.24483, 48.93617, 47.23159,
    41.8115, 40.59438,
  46.67609, 47.29061, 47.90333, 48.5539, 49.21495, 50.08963, 50.36596,
    50.24707, 50.57861, 51.12508, 51.34843, 51.74409, 51.49311, 50.4459,
    51.06807, 51.72923, 50.55424, 49.42, 50.35038, 51.47914, 54.13725,
    55.11119, 53.06168, 57.99381, 60.07177, 52.91412, 51.77975, 46.34397,
    41.77022, 39.6556,
  52.30434, 52.70984, 53.49564, 54.33269, 54.86239, 55.14342, 55.31631,
    55.47325, 56.24869, 56.8505, 56.68802, 56.76663, 56.45049, 56.00046,
    55.32589, 54.79068, 53.35074, 51.59898, 51.79882, 56.74335, 58.51825,
    50.89537, 50.92527, 52.53147, 54.46456, 53.14663, 49.16608, 48.89711,
    47.95832, 41.84294,
  56.745, 57.8339, 59.09066, 60.64368, 60.65556, 60.19257, 60.83555,
    61.22528, 61.20817, 61.91644, 62.81242, 65.05521, 67.13696, 65.53725,
    63.34231, 67.54707, 68.48047, 64.33552, 54.41898, 55.04858, 52.3971,
    49.06995, 49.89343, 51.1391, 53.52832, 52.03079, 54.37926, 64.96931,
    60.45527, 40.64093,
  61.91441, 63.68597, 65.36287, 67.20447, 67.95071, 68.57203, 69.28837,
    69.42097, 68.93318, 68.63575, 68.45924, 67.9509, 64.52762, 63.08046,
    66.3748, 67.4325, 64.63263, 55.86377, 52.23758, 51.62709, 50.01172,
    49.13682, 49.8119, 52.21751, 53.00595, 49.25419, 58.33737, 65.61249,
    58.15086, 38.86367,
  67.77497, 69.04942, 69.32729, 69.51373, 69.12702, 69.01309, 69.47147,
    69.22937, 66.46659, 65.07077, 63.22476, 61.01583, 58.70338, 57.29575,
    56.51536, 55.76843, 54.52303, 52.93705, 50.03306, 49.47454, 48.59345,
    48.44917, 50.0774, 52.09459, 50.8533, 48.47583, 59.62278, 64.35965,
    45.64771, 39.53032,
  69.23969, 69.51576, 69.65652, 69.57296, 69.0929, 68.98172, 67.71812,
    65.00777, 64.58321, 63.7285, 62.58294, 61.40886, 60.36058, 62.90753,
    63.66829, 56.78547, 55.29045, 56.43156, 55.62886, 52.2716, 49.95534,
    52.25581, 56.68855, 56.59084, 51.64472, 51.80783, 54.73462, 51.22225,
    41.79056, 39.41944,
  71.02675, 71.60976, 71.75084, 71.90765, 71.30163, 70.00196, 65.34479,
    66.58698, 67.01113, 68.61085, 70.58739, 71.02799, 70.77618, 68.23658,
    63.07534, 62.64418, 62.59871, 61.44117, 58.83679, 57.42171, 57.92548,
    57.29881, 56.25922, 52.23044, 59.41684, 67.39735, 58.11645, 42.31543,
    39.64341, 38.39686,
  74.47282, 74.55982, 74.80184, 74.09428, 73.82195, 73.47307, 72.80029,
    72.90356, 73.24531, 75.25015, 76.58227, 70.56189, 66.28135, 63.93233,
    61.97695, 61.02909, 60.80593, 59.54732, 57.68979, 56.61723, 58.18692,
    55.96575, 50.44113, 46.64087, 48.46645, 49.89008, 43.84885, 39.22633,
    38.86456, 38.28009,
  80.06509, 76.6297, 79.85746, 80.99419, 80.54359, 79.02376, 77.91666,
    74.73648, 71.62153, 72.1217, 71.51795, 68.46069, 69.19181, 68.0664,
    61.17918, 59.48092, 56.8553, 55.20707, 53.46128, 52.66203, 53.98793,
    51.59578, 45.43868, 49.79544, 52.21672, 42.06855, 39.01245, 39.39692,
    39.14288, 38.57498,
  86.7722, 87.40551, 90.18072, 90.40342, 88.84613, 84.52203, 76.65704,
    72.27091, 72.33982, 70.67371, 70.75624, 69.84613, 69.65998, 69.44281,
    63.75499, 57.61032, 55.26714, 53.26195, 51.5528, 52.61065, 52.54886,
    48.3111, 44.75874, 48.21318, 49.78043, 41.10094, 39.53139, 39.70657,
    39.81417, 38.98021,
  84.41366, 86.82095, 85.8284, 82.90231, 79.97979, 78.11157, 77.50684,
    77.20936, 74.47772, 73.59406, 74.72924, 73.26397, 73.96312, 73.45074,
    70.59021, 67.90742, 56.09646, 57.00988, 57.00484, 56.00584, 50.97779,
    49.88029, 52.82257, 44.91875, 41.44128, 40.42748, 39.55297, 39.16015,
    39.37919, 38.9021,
  75.9785, 75.63501, 74.52725, 73.18373, 72.09515, 73.86309, 79.18318,
    78.99436, 75.63254, 74.95033, 74.02716, 72.33131, 70.78078, 70.67752,
    69.85774, 62.5944, 60.41208, 57.89693, 58.51104, 59.68082, 55.29337,
    48.70008, 43.36878, 41.17919, 40.31534, 40.33508, 39.55893, 39.01758,
    38.81963, 38.53816,
  72.2647, 72.40607, 72.57303, 72.2792, 72.07014, 72.87639, 73.68417,
    73.31992, 72.51012, 71.56982, 71.1667, 70.04799, 68.9892, 68.61906,
    64.37219, 59.62343, 57.74255, 53.76793, 52.53356, 50.88229, 44.76884,
    42.90823, 40.88706, 40.43143, 40.48588, 40.25452, 39.56828, 39.06704,
    38.78951, 38.4795,
  71.47207, 71.67815, 71.66531, 71.58281, 71.7483, 71.2187, 71.24517,
    71.79507, 71.44051, 70.77435, 69.53511, 69.3364, 69.80363, 66.8476,
    60.56271, 56.43287, 52.97506, 49.93333, 50.96846, 49.91778, 42.31053,
    42.51233, 41.41331, 40.49483, 40.11861, 40.15381, 39.47496, 38.76382,
    38.61718, 38.45223,
  70.55381, 71.09484, 70.78295, 70.7674, 70.41171, 70.26292, 70.05582,
    70.26208, 70.60252, 69.84189, 69.61755, 69.85611, 68.50774, 64.5811,
    62.31004, 55.79869, 49.68861, 46.86691, 49.39341, 48.2851, 42.70169,
    42.48525, 41.46254, 40.61359, 39.69054, 39.57745, 39.22197, 38.57638,
    38.44863, 38.33879,
  71.93204, 71.73719, 70.53381, 69.6641, 69.74505, 69.32115, 69.01273,
    68.90212, 67.62018, 66.50082, 67.55998, 65.02496, 58.35828, 56.77922,
    54.98476, 52.49881, 52.46979, 53.21872, 55.74297, 54.56026, 48.03465,
    43.80119, 41.42186, 40.70969, 39.48166, 39.14915, 38.96156, 38.56644,
    38.4028, 38.32751,
  71.93065, 71.41576, 68.96447, 66.43497, 65.73499, 65.03767, 64.42388,
    63.77128, 63.18056, 64.62527, 64.15462, 58.7268, 56.05387, 54.36492,
    52.54794, 51.20642, 52.06318, 53.44366, 54.31863, 54.1532, 50.44021,
    45.50563, 41.78103, 40.95779, 39.90554, 39.21751, 38.92959, 38.59491,
    38.39653, 38.33415,
  69.932, 68.28865, 65.38087, 63.1117, 62.20259, 61.65042, 61.15265,
    60.76206, 61.12179, 62.52821, 60.55802, 56.67388, 56.19489, 54.55881,
    52.18016, 49.94624, 49.09472, 48.66359, 48.79134, 48.18358, 46.95804,
    46.02721, 43.91641, 41.93111, 40.51329, 39.59193, 38.95435, 38.62242,
    38.41662, 38.32875,
  69.05092, 66.0968, 63.6364, 61.99134, 61.23426, 60.20249, 60.02622,
    59.82372, 61.22121, 61.68633, 58.30057, 55.60325, 54.45473, 51.92343,
    49.12763, 47.3448, 46.05554, 45.22197, 44.88384, 44.1909, 45.5703,
    46.57093, 44.64976, 44.90595, 42.637, 40.30285, 39.12722, 38.81842,
    38.48658, 38.34151,
  67.7494, 65.95663, 63.22481, 61.8146, 62.19748, 62.21914, 61.26503,
    59.73346, 59.99616, 58.74296, 55.06753, 53.36094, 51.55341, 49.21618,
    46.77488, 45.85926, 45.39203, 44.02743, 43.29648, 42.92302, 44.25288,
    45.02494, 42.72594, 43.8075, 43.99935, 41.65592, 39.65672, 39.42844,
    38.86421, 38.39338,
  68.14867, 66.91389, 65.50754, 64.64954, 63.96999, 62.99913, 62.67934,
    61.84113, 61.60486, 57.99196, 53.8462, 53.10851, 51.64339, 49.91164,
    47.96191, 46.75886, 46.31955, 45.1808, 43.61155, 42.99521, 43.13915,
    43.05815, 42.37469, 42.1974, 42.91344, 43.24815, 41.48162, 39.93698,
    39.31158, 38.59206,
  68.07915, 68.50848, 65.06307, 63.4113, 63.08514, 62.11515, 60.79663,
    60.22375, 61.09269, 58.27551, 53.8451, 53.54387, 52.42479, 50.54211,
    48.60748, 47.6098, 46.63136, 45.93246, 44.67414, 43.23296, 43.11965,
    43.15536, 42.73921, 41.99707, 41.42942, 42.53978, 42.73831, 41.1091,
    40.27674, 39.22081,
  68.9824, 70.69217, 68.48898, 65.26401, 63.08966, 61.6114, 62.05247,
    62.62989, 60.71497, 57.49982, 55.35773, 54.797, 53.62639, 50.79202,
    48.04745, 46.9994, 46.36753, 46.01615, 45.2212, 43.74042, 43.63791,
    43.68274, 42.53237, 41.56076, 41.45775, 41.90812, 42.91231, 42.055,
    40.17288, 39.06673,
  69.83642, 70.47938, 66.94068, 64.32154, 63.00842, 61.47382, 62.09469,
    61.88811, 58.80014, 56.44768, 55.92471, 55.06816, 53.14006, 50.27707,
    47.96561, 46.67242, 45.96866, 45.82235, 45.10457, 43.90034, 44.47738,
    46.08571, 46.26209, 44.65129, 43.77739, 43.71215, 44.75616, 44.21977,
    40.44181, 38.45132,
  69.33284, 68.53419, 66.14732, 65.28204, 64.77937, 63.31456, 62.62512,
    60.43943, 56.75032, 55.98715, 55.32729, 54.33224, 52.37268, 49.93144,
    48.59091, 47.50199, 46.51044, 46.54546, 46.85569, 47.08273, 47.81701,
    47.92586, 46.63047, 45.31562, 44.6132, 44.53461, 44.3359, 45.66158,
    43.99218, 39.53559,
  66.73479, 65.59891, 65.94312, 66.56815, 66.22144, 66.0764, 63.56075,
    58.44804, 55.77467, 55.50193, 54.25308, 52.90034, 51.37786, 50.31549,
    50.17233, 49.98062, 49.84168, 50.0401, 48.86372, 47.045, 46.44143,
    45.65242, 44.3493, 43.44424, 43.37601, 43.53611, 43.23019, 42.48288,
    42.42523, 40.30965,
  65.59045, 65.39318, 64.89021, 63.81708, 63.56138, 65.24714, 64.99113,
    59.75805, 56.69502, 57.44914, 57.67025, 57.24364, 55.78212, 54.26011,
    52.98706, 51.70189, 49.68222, 47.47819, 46.20498, 44.66625, 43.52956,
    43.0019, 42.51185, 42.11023, 41.84264, 41.93322, 41.62672, 40.63184,
    39.63061, 38.60666,
  33.02636, 33.06883, 33.11969, 33.16751, 33.16242, 33.17242, 33.20924,
    33.2758, 33.39219, 33.55224, 34.44285, 34.62243, 33.40468, 33.52243,
    33.66061, 33.33882, 33.25513, 33.35482, 33.43758, 34.0402, 34.37188,
    33.84062, 33.93113, 34.65636, 35.13899, 34.88813, 37.18357, 38.65747,
    34.95919, 33.67333,
  33.67009, 33.78664, 33.60139, 33.88712, 33.73347, 33.61745, 33.73795,
    33.8532, 33.98558, 34.17403, 34.54346, 35.08619, 35.41151, 34.67424,
    34.24392, 34.38562, 33.87772, 34.05976, 34.63381, 35.24666, 35.30696,
    35.00779, 35.38148, 36.42583, 40.98821, 42.55443, 37.64623, 40.02824,
    35.54155, 34.10648,
  33.93577, 34.00856, 33.99753, 34.05908, 34.07595, 34.12618, 34.16303,
    34.27818, 34.41793, 34.51673, 34.6811, 35.08496, 35.37887, 35.83902,
    36.11983, 35.43476, 35.48311, 36.10981, 36.43882, 37.04254, 38.35107,
    40.01595, 41.12469, 40.59724, 45.17266, 48.31813, 40.01171, 39.47067,
    35.54557, 34.7294,
  34.93274, 35.09207, 35.37765, 35.67052, 36.00578, 36.58598, 36.70617,
    36.48169, 36.61924, 36.97281, 37.06698, 37.33992, 37.26241, 36.85985,
    38.00462, 39.21345, 38.75381, 37.99408, 38.70731, 39.60822, 41.95865,
    43.17326, 41.60832, 46.54652, 49.26123, 43.02413, 42.51429, 38.7779,
    35.50911, 34.03543,
  37.28685, 37.33128, 37.7908, 38.31644, 38.63404, 38.78855, 38.82872,
    38.81168, 39.38938, 39.77031, 39.43081, 39.42465, 39.39763, 39.67857,
    40.32124, 41.0157, 40.49087, 39.86725, 40.36086, 45.18662, 47.22543,
    40.48082, 40.42006, 41.92239, 43.68914, 42.63654, 39.89074, 39.63046,
    39.68576, 35.72403,
  39.73075, 40.31752, 41.19272, 42.27637, 42.14097, 41.61337, 41.90993,
    42.05886, 41.97365, 42.36354, 42.79082, 44.48587, 46.45219, 46.29818,
    45.25433, 53.86936, 64.2597, 51.7421, 43.11317, 44.26527, 42.31009,
    39.12265, 39.55922, 40.31171, 42.34724, 41.41768, 44.39512, 58.7983,
    52.58907, 34.83789,
  42.51461, 43.46442, 44.56989, 45.8102, 46.19201, 46.53456, 47.92679,
    49.82539, 50.31847, 50.26179, 50.4734, 49.30437, 47.17963, 46.44098,
    51.82979, 59.88279, 54.40332, 45.12751, 41.95535, 41.4245, 39.9659,
    39.10862, 39.57274, 41.41393, 42.41307, 39.29833, 49.09439, 66.7584,
    51.79016, 33.37433,
  46.07203, 47.52721, 49.11535, 50.77403, 51.05453, 52.94336, 55.07784,
    52.75736, 50.57304, 50.06308, 48.83891, 46.82162, 44.72907, 43.73447,
    44.27826, 45.01289, 43.8107, 42.44016, 40.33587, 39.8786, 39.13852,
    38.84993, 40.07434, 41.72125, 41.09107, 38.80985, 50.88301, 57.65815,
    39.25082, 34.32985,
  51.86448, 53.01471, 54.20729, 54.5607, 54.08279, 54.66623, 52.86739,
    50.98082, 50.52875, 49.60435, 48.0337, 46.21061, 44.76883, 46.903,
    48.15552, 43.60267, 43.22116, 44.5491, 44.05166, 41.49304, 39.47785,
    40.94917, 44.56514, 44.82932, 41.01155, 41.31653, 45.35225, 44.07032,
    36.54668, 34.25884,
  58.06219, 60.27919, 60.7188, 60.97108, 59.0303, 54.53949, 49.66703,
    49.80023, 49.39878, 49.58175, 50.45784, 53.14187, 52.92113, 49.97093,
    46.67419, 46.75117, 47.40041, 46.99647, 45.40897, 44.84223, 45.30987,
    45.44459, 45.61197, 43.07801, 49.40745, 60.51287, 49.82313, 36.9142,
    34.56533, 33.173,
  68.69952, 68.24462, 68.24022, 65.75508, 63.63699, 60.64035, 56.7107,
    58.85476, 60.37494, 69.53494, 71.6188, 53.75822, 47.38376, 45.76347,
    44.79126, 44.88529, 45.91657, 46.56432, 45.12043, 44.61445, 47.1283,
    46.2252, 41.98476, 39.00895, 41.88497, 44.55519, 38.83644, 34.0942,
    33.59701, 33.02148,
  72.7921, 68.42421, 71.29597, 72.24345, 72.69724, 71.70615, 71.58272,
    69.59441, 58.9655, 61.9654, 60.73207, 47.50585, 48.82512, 49.02922,
    44.3772, 45.29824, 44.2177, 43.73824, 42.70024, 42.68162, 45.23193,
    43.58183, 38.14349, 41.80948, 44.09018, 36.3345, 33.63964, 34.0541,
    33.86119, 33.27959,
  76.50001, 76.87859, 81.82929, 82.53931, 82.73939, 79.82615, 72.16052,
    61.40838, 61.59846, 57.09217, 55.70707, 49.66358, 52.81364, 53.36799,
    45.93731, 44.87186, 44.30925, 42.9348, 41.62668, 43.47491, 44.59127,
    40.70247, 37.44921, 41.73406, 43.45713, 35.42038, 33.9781, 34.23347,
    34.44138, 33.64614,
  78.13972, 83.51952, 82.06022, 79.51151, 76.58131, 73.43089, 70.85733,
    70.39459, 69.03507, 68.1596, 69.65966, 69.75263, 71.90874, 73.03059,
    65.89199, 52.9147, 44.31987, 45.84497, 46.93869, 47.35235, 43.39074,
    42.04926, 44.47467, 38.78397, 36.02044, 34.72979, 33.97585, 33.7046,
    34.03735, 33.58001,
  72.15508, 72.20964, 70.72162, 69.02695, 67.37171, 68.30869, 73.16055,
    73.43028, 70.85999, 70.39748, 70.13637, 68.98045, 55.95983, 61.15621,
    65.02621, 48.41467, 48.19299, 47.51008, 50.60953, 52.27653, 46.75161,
    42.03247, 37.74119, 35.37856, 34.49686, 34.7621, 34.05757, 33.58636,
    33.50275, 33.25225,
  68.56652, 67.29461, 66.42199, 65.57011, 66.19905, 67.1416, 68.12412,
    67.96161, 67.57651, 64.19907, 59.4014, 52.76758, 49.4632, 51.62537,
    50.21181, 47.24476, 47.72482, 45.34245, 45.73266, 45.23134, 39.09743,
    36.71052, 34.75399, 34.58971, 34.87325, 34.72752, 34.15393, 33.67621,
    33.45199, 33.18156,
  64.8916, 63.23674, 62.3334, 62.03462, 62.26596, 61.48503, 60.43849,
    59.72621, 57.9333, 55.42632, 51.04123, 51.2549, 54.67203, 51.15452,
    47.72607, 46.25727, 44.53659, 42.2206, 44.10904, 43.45044, 35.79359,
    35.97385, 35.32083, 34.72919, 34.58653, 34.67361, 34.0835, 33.42132,
    33.30917, 33.15892,
  60.64796, 60.14476, 58.85679, 58.23209, 57.21637, 56.51929, 55.94564,
    55.42236, 54.42075, 52.16074, 51.73916, 53.59413, 51.70639, 50.37729,
    51.27137, 47.29219, 42.07885, 39.28036, 42.52191, 42.02739, 36.24673,
    36.3317, 35.77611, 35.13116, 34.1739, 34.16473, 33.83719, 33.22793,
    33.14, 33.05979,
  59.83572, 58.62725, 55.89201, 53.99725, 53.29394, 52.47086, 52.11568,
    52.04483, 50.96325, 49.90017, 51.19905, 49.55925, 43.98829, 43.97382,
    44.35017, 43.02747, 43.12465, 43.70324, 46.77414, 46.22462, 40.26931,
    37.43879, 36.0756, 35.32443, 34.05196, 33.79299, 33.61126, 33.2276,
    33.09939, 33.02668,
  57.40924, 55.87743, 53.31575, 51.28046, 50.7786, 50.28866, 49.90002,
    49.42865, 48.79263, 50.03809, 49.56373, 43.90216, 41.01498, 40.62291,
    40.35258, 39.83351, 41.28693, 43.29755, 45.36737, 46.31919, 43.23996,
    39.22908, 36.32029, 35.47378, 34.49788, 33.87627, 33.57708, 33.27905,
    33.10696, 33.03505,
  54.50024, 53.5797, 51.69874, 49.70715, 48.96297, 48.46475, 47.8885,
    47.23929, 47.16208, 48.20555, 45.35404, 40.43444, 40.36332, 40.52259,
    40.18378, 39.29916, 39.30408, 39.57773, 40.67642, 41.10353, 40.43172,
    39.85104, 38.26319, 36.30235, 34.99552, 34.2301, 33.60384, 33.2846,
    33.12617, 33.04702,
  53.52227, 52.17918, 50.10117, 48.5586, 47.71213, 46.58373, 46.09428,
    45.54964, 46.6852, 46.86211, 42.75189, 39.77337, 39.96344, 39.78818,
    39.18569, 38.60025, 37.92464, 37.46314, 37.44387, 37.07152, 38.6524,
    39.76734, 39.04028, 39.62676, 37.38818, 34.98311, 33.77909, 33.48766,
    33.1772, 33.05257,
  52.43934, 50.90895, 48.39121, 46.97183, 47.27439, 47.4127, 46.81258,
    45.72519, 46.49148, 45.27618, 41.04946, 39.50829, 39.10818, 38.80854,
    38.09028, 38.05349, 37.87646, 36.68249, 36.07139, 35.93441, 37.52308,
    38.21967, 36.79557, 38.46014, 38.86702, 36.29233, 34.20471, 34.05962,
    33.56239, 33.12578,
  51.40914, 49.91139, 48.87873, 48.34363, 48.21132, 48.11734, 48.64951,
    48.72109, 49.35773, 45.74146, 40.67847, 39.84206, 39.48585, 39.53017,
    39.12354, 38.74197, 38.7561, 37.82432, 36.42885, 36.08968, 36.56062,
    36.6339, 36.11882, 36.32502, 37.49279, 37.83259, 35.97353, 34.51315,
    33.966, 33.30615,
  50.86628, 51.56208, 48.90717, 47.94804, 48.29758, 48.2063, 47.84141,
    48.01412, 49.34573, 45.91728, 40.49219, 39.87205, 39.79658, 39.66277,
    39.40138, 39.42828, 38.97542, 38.67586, 37.49738, 36.0624, 36.35033,
    36.71999, 36.50347, 35.80721, 35.26742, 36.54976, 36.84767, 35.41775,
    34.87314, 33.86976,
  52.03703, 54.05689, 52.63203, 50.34252, 48.70862, 47.62288, 48.66228,
    49.95479, 48.36701, 44.44321, 41.17365, 40.51584, 40.58173, 39.79124,
    38.83902, 38.80008, 38.6444, 38.67377, 37.99345, 36.48655, 36.84431,
    37.23195, 36.07911, 35.1906, 35.05733, 35.61034, 36.96568, 36.30843,
    34.75826, 33.72027,
  53.30485, 54.42572, 51.25826, 49.16247, 48.12284, 47.02805, 48.39939,
    49.07027, 45.90329, 42.79579, 41.45654, 40.77705, 40.25694, 39.37355,
    38.84954, 38.50914, 38.24048, 38.46892, 37.83072, 36.43605, 37.22527,
    39.19112, 39.47888, 37.80289, 36.94609, 37.09217, 38.61347, 38.45035,
    34.98495, 33.12453,
  52.51019, 52.05476, 49.959, 49.34201, 49.41927, 48.72477, 49.09556,
    47.50544, 43.64901, 42.35093, 41.148, 40.37363, 39.80191, 39.20327,
    39.42888, 39.12927, 38.32246, 38.45413, 38.64589, 38.57077, 39.97643,
    40.9583, 39.83216, 38.27761, 37.53119, 37.67749, 37.79113, 39.6381,
    38.21393, 34.09505,
  49.75862, 48.64394, 49.11935, 50.41448, 51.1631, 52.10368, 50.5476,
    46.08537, 43.19799, 42.32257, 40.30234, 38.74192, 38.03878, 38.50585,
    39.8366, 40.34401, 40.50742, 41.20764, 40.17123, 38.44778, 38.47237,
    38.12945, 36.96629, 36.17799, 36.27911, 36.68916, 36.68135, 36.41222,
    36.8321, 34.80527,
  48.84029, 48.84518, 48.68527, 48.23452, 48.57097, 51.13911, 51.78095,
    46.69524, 43.20169, 43.09688, 42.34693, 41.63725, 41.10647, 41.65009,
    42.38238, 42.16672, 40.98164, 39.43745, 38.27944, 36.89272, 36.0819,
    35.74073, 35.48259, 35.28599, 35.26384, 35.66496, 35.68545, 34.95532,
    34.20712, 33.32852,
  23.71678, 23.76854, 23.80622, 23.84324, 23.83076, 23.82301, 23.84658,
    23.88153, 23.94448, 24.08622, 25.05237, 25.21221, 24.06777, 24.19527,
    24.34865, 23.9914, 23.85891, 23.93232, 23.96853, 24.55544, 24.87388,
    24.3322, 24.36144, 24.98401, 25.3494, 25.04231, 27.60794, 29.43835,
    25.84898, 24.47773,
  24.15661, 24.24746, 24.04833, 24.33681, 24.17272, 24.01614, 24.09248,
    24.17366, 24.28329, 24.48356, 24.93112, 25.54357, 25.88495, 25.09598,
    24.66593, 24.73994, 24.17162, 24.25319, 24.75771, 25.31662, 25.29355,
    24.84355, 24.99583, 25.94416, 30.32813, 31.35156, 28.12269, 31.30952,
    26.60254, 25.07459,
  24.15664, 24.19502, 24.1869, 24.24554, 24.22715, 24.22638, 24.24957,
    24.33261, 24.44123, 24.51999, 24.65654, 25.08874, 25.38497, 25.80673,
    25.96096, 25.14806, 25.07122, 25.50749, 25.59637, 25.94792, 26.90074,
    28.33401, 29.39854, 29.11714, 34.00134, 36.87238, 30.56876, 30.79813,
    26.53414, 25.70801,
  24.45566, 24.52461, 24.74976, 24.95059, 25.24163, 25.80723, 25.8982,
    25.61504, 25.67284, 26.02894, 26.15324, 26.38666, 26.15573, 25.71564,
    26.80086, 27.92103, 27.32273, 26.25499, 26.59948, 27.19112, 29.58255,
    30.91282, 29.85336, 34.56902, 36.8709, 32.86164, 33.38501, 30.19735,
    26.55012, 24.91658,
  25.72163, 25.58301, 25.92756, 26.31502, 26.64712, 26.82622, 26.77416,
    26.64712, 27.20373, 27.64312, 27.35479, 27.18688, 26.93102, 27.21312,
    28.01107, 28.71078, 28.00687, 27.18601, 27.76254, 32.28293, 34.00634,
    28.80421, 28.72479, 30.59499, 32.61324, 32.20682, 30.39005, 30.698,
    31.27755, 26.80279,
  27.21576, 27.49636, 28.27325, 29.34083, 29.24521, 28.66831, 28.70887,
    28.58771, 28.21197, 28.25242, 28.26744, 29.8618, 31.95622, 32.03716,
    31.51792, 39.34072, 47.62727, 37.6883, 31.02282, 32.60033, 30.78981,
    27.49644, 27.91509, 28.80869, 31.4047, 30.94145, 33.72445, 46.95179,
    42.30311, 26.09935,
  29.41865, 29.94179, 30.76602, 31.80095, 31.99973, 31.9248, 32.88714,
    34.56194, 34.78594, 34.4721, 34.62879, 33.65481, 31.99991, 32.0676,
    37.6228, 45.47144, 42.08035, 33.43293, 30.4216, 29.9914, 28.398,
    27.42077, 27.87264, 30.15376, 31.67394, 29.10972, 38.77229, 54.80732,
    41.68091, 24.52743,
  31.99001, 32.79734, 33.96413, 35.2711, 35.41114, 37.59247, 40.13025,
    37.97091, 35.92488, 35.35544, 34.19173, 32.27401, 30.50805, 30.26491,
    31.97799, 33.48183, 32.39116, 30.89291, 28.83227, 28.40616, 27.6375,
    27.27093, 28.53319, 30.86202, 30.5936, 28.84581, 41.11457, 47.20827,
    30.75652, 24.81386,
  36.37734, 37.17918, 38.48783, 39.05207, 39.22264, 40.89382, 39.867,
    38.03593, 37.53197, 36.43473, 34.39365, 32.14281, 30.58218, 33.52147,
    35.57151, 31.38427, 31.05911, 32.74038, 32.69674, 30.09845, 27.69794,
    29.15727, 33.29696, 34.17738, 30.62035, 31.04894, 36.89463, 35.52814,
    26.92517, 24.84248,
  42.08245, 44.59632, 46.24624, 47.90608, 47.09908, 42.85439, 38.17031,
    37.87448, 36.77003, 35.58198, 35.44742, 38.00674, 38.4343, 36.36725,
    33.84472, 33.89595, 34.83323, 35.3408, 33.56432, 31.71471, 31.96599,
    32.41348, 33.12987, 31.2993, 37.01979, 47.69079, 39.46992, 27.57478,
    25.26707, 23.97259,
  58.73119, 61.35275, 56.2549, 50.09378, 48.07657, 46.60817, 42.49906,
    44.08958, 45.53042, 53.10435, 57.28904, 39.21032, 33.29309, 31.9241,
    31.13238, 31.98304, 33.15145, 33.03417, 31.84206, 31.56163, 34.12497,
    33.41436, 30.24568, 28.01064, 31.447, 35.26041, 29.84367, 24.69578,
    24.37094, 23.79938,
  74.28508, 61.38707, 65.99919, 68.23263, 66.56519, 56.77492, 58.34174,
    54.09509, 45.59734, 49.12571, 47.54464, 32.71858, 33.22153, 33.78574,
    30.98591, 31.43904, 30.77151, 30.48423, 30.06267, 30.68494, 33.4367,
    32.06028, 27.63569, 31.08631, 33.00404, 26.6936, 24.38938, 24.76249,
    24.60819, 24.0169,
  74.1581, 73.88833, 78.43401, 80.51269, 82.46169, 81.32652, 70.13583,
    48.05139, 46.691, 42.95926, 39.34538, 32.33082, 36.47364, 38.19584,
    32.61976, 31.34933, 31.1618, 30.35516, 29.75975, 31.94333, 33.47786,
    30.05042, 27.11547, 31.84435, 33.37714, 25.94777, 24.57676, 24.89103,
    25.13446, 24.33816,
  76.30253, 81.81801, 82.48368, 81.41906, 79.81982, 75.96481, 73.71575,
    69.83978, 59.64833, 55.40998, 61.99773, 59.54156, 60.01313, 57.48626,
    48.81988, 38.35272, 31.483, 33.37034, 34.9075, 35.86631, 32.53643,
    31.26202, 33.22318, 29.21495, 26.72477, 25.1912, 24.56883, 24.37034,
    24.74677, 24.27238,
  67.36699, 71.4325, 66.42594, 61.51566, 55.56146, 63.92392, 74.56009,
    75.37686, 73.25905, 72.95373, 71.65754, 54.72446, 42.59272, 47.51535,
    49.43331, 35.21612, 35.248, 35.34457, 38.2695, 39.41669, 35.45096,
    31.65886, 28.50137, 25.99601, 24.89906, 25.21256, 24.61667, 24.25163,
    24.23268, 23.98135,
  53.59624, 51.72028, 50.3036, 48.84802, 49.21783, 54.70249, 61.03661,
    59.30801, 56.3229, 53.15281, 48.1532, 39.53759, 34.48704, 37.4172,
    36.83543, 34.60222, 35.81559, 34.19703, 35.08391, 34.79544, 29.6134,
    27.07533, 25.19319, 25.12362, 25.41309, 25.18037, 24.71048, 24.36348,
    24.21084, 23.93274,
  48.93563, 47.02853, 46.10385, 46.19595, 47.3707, 48.09726, 48.26641,
    47.9897, 46.09043, 42.88301, 37.41221, 35.80558, 38.85169, 36.97211,
    35.06925, 34.59685, 33.63798, 31.83838, 33.72023, 32.76527, 25.91298,
    26.03553, 25.71687, 25.31287, 25.17437, 25.19443, 24.65971, 24.13483,
    24.08006, 23.89516,
  44.99073, 44.92493, 44.60218, 45.12363, 45.13165, 45.38371, 45.11556,
    44.35135, 42.87106, 38.88063, 37.06534, 38.69617, 38.32623, 37.77341,
    39.33555, 36.34068, 31.71659, 29.2297, 32.3547, 31.59418, 26.29436,
    26.53934, 26.21376, 25.64281, 24.75018, 24.79045, 24.48107, 23.94636,
    23.89705, 23.80712,
  46.02695, 46.25657, 44.51929, 43.43005, 43.09798, 42.45302, 41.96483,
    41.32949, 39.48987, 37.09256, 37.70366, 36.77745, 32.41388, 32.86411,
    33.69983, 32.41857, 32.06123, 32.50131, 35.45144, 34.70362, 29.50937,
    27.46158, 26.52233, 25.80008, 24.66096, 24.44711, 24.29379, 23.94199,
    23.84588, 23.78335,
  46.48016, 46.03955, 43.76733, 41.70121, 41.21539, 40.74298, 40.3046,
    39.57306, 38.13931, 38.24521, 37.53078, 32.52213, 29.63481, 29.48907,
    29.26138, 28.68766, 30.10362, 32.15822, 34.417, 35.26715, 32.5511,
    29.24618, 26.77293, 25.93042, 25.04679, 24.50364, 24.25687, 23.9857,
    23.84573, 23.78465,
  45.22202, 44.58089, 42.41228, 40.6421, 40.07286, 39.84917, 39.47981,
    38.61115, 37.77693, 37.93711, 34.4242, 29.04861, 28.70179, 28.91689,
    28.61269, 27.9602, 28.22741, 28.82384, 30.25406, 30.99756, 30.57537,
    30.05073, 28.57635, 26.67398, 25.42718, 24.76525, 24.25938, 23.98167,
    23.86073, 23.78714,
  45.08302, 43.32628, 41.5906, 40.3513, 39.8372, 39.05532, 38.62873,
    37.65446, 37.59342, 36.38123, 31.21096, 27.80103, 28.09958, 28.22478,
    27.98641, 27.69621, 27.33075, 27.19276, 27.39483, 27.27176, 28.57495,
    29.28792, 29.16081, 29.62113, 27.63437, 25.38807, 24.38836, 24.13441,
    23.89476, 23.80001,
  43.96082, 42.8671, 40.7902, 39.49725, 39.79425, 39.94292, 39.09391,
    37.47977, 37.04357, 34.27922, 29.20509, 27.56346, 27.61395, 27.72736,
    27.37152, 27.63725, 27.59307, 26.59582, 26.13474, 26.0952, 27.45543,
    27.85607, 27.13362, 28.84621, 29.07407, 26.48762, 24.73154, 24.61354,
    24.19284, 23.83267,
  43.05487, 41.98901, 40.87938, 40.29788, 40.22414, 40.14962, 40.31904,
    39.71661, 39.13281, 34.36491, 28.94173, 28.19831, 28.3077, 28.70818,
    28.5464, 28.41258, 28.4857, 27.59174, 26.42079, 26.27543, 26.76385,
    26.76668, 26.45308, 26.79357, 27.96768, 28.10642, 26.30645, 24.98449,
    24.54197, 23.96847,
  42.17036, 42.76752, 40.33735, 39.51051, 39.87515, 39.81572, 39.44682,
    39.2787, 39.53299, 34.80761, 29.07328, 28.48233, 28.72088, 28.919,
    28.93836, 29.02498, 28.69906, 28.46001, 27.32355, 26.15694, 26.53285,
    26.84377, 26.68144, 26.00774, 25.67798, 27.02379, 27.16805, 25.7909,
    25.42376, 24.42536,
  42.05494, 43.9866, 42.89731, 41.29488, 39.97714, 39.16573, 40.20444,
    41.12345, 38.74315, 33.62666, 29.68013, 29.00596, 29.34185, 28.91169,
    28.34751, 28.45843, 28.35407, 28.48947, 27.7743, 26.43946, 26.97013,
    27.25137, 26.19648, 25.42632, 25.29609, 25.97158, 27.37547, 26.61748,
    25.43839, 24.3728,
  42.91665, 44.1823, 42.001, 40.43537, 39.60578, 38.90799, 40.28244,
    40.58614, 36.48175, 31.99018, 29.81404, 29.16054, 29.05236, 28.59204,
    28.28679, 28.10315, 28.00275, 28.33171, 27.64532, 26.34068, 27.15312,
    28.8173, 28.92439, 27.529, 26.90501, 27.10678, 28.91366, 28.62178,
    25.47415, 23.84456,
  42.78307, 42.90555, 41.13689, 40.6173, 41.01273, 40.67528, 41.10417,
    39.01634, 34.09066, 31.30038, 29.42315, 28.79958, 28.69545, 28.52156,
    28.8844, 28.63956, 27.96681, 28.08797, 28.18074, 28.00316, 29.39807,
    30.17288, 29.1956, 27.83536, 27.39389, 27.60868, 28.02972, 30.03666,
    28.45495, 24.63679,
  40.46281, 39.7777, 40.30632, 41.59563, 42.71714, 44.05426, 42.59362,
    37.76083, 33.70781, 31.40484, 28.70404, 27.28165, 27.05023, 27.75879,
    29.02312, 29.43039, 29.5099, 30.10562, 29.18601, 27.81456, 27.96552,
    27.64821, 26.60205, 25.98543, 26.22, 26.77909, 26.91808, 26.94022,
    27.52707, 25.26363,
  39.28175, 39.51154, 39.56889, 39.39736, 39.97015, 42.86887, 43.46532,
    37.86327, 33.32026, 31.68034, 30.14687, 29.45866, 29.38567, 30.25212,
    31.03992, 30.9577, 29.88648, 28.53512, 27.55735, 26.38309, 25.74319,
    25.53742, 25.34686, 25.28423, 25.3954, 25.93889, 26.11624, 25.47909,
    24.88905, 24.05807,
  17.21845, 17.24786, 17.27626, 17.30108, 17.28836, 17.28526, 17.30391,
    17.32797, 17.37545, 17.44251, 18.21923, 18.33761, 17.46813, 17.60441,
    17.73426, 17.43442, 17.32892, 17.36065, 17.37738, 17.86694, 18.10322,
    17.64251, 17.62224, 18.1039, 18.36679, 18.04801, 20.26277, 21.81756,
    19.06623, 17.89275,
  17.51968, 17.56397, 17.40266, 17.62378, 17.5013, 17.371, 17.41702,
    17.48078, 17.5563, 17.70706, 18.06279, 18.604, 18.91337, 18.24807,
    17.93906, 17.96558, 17.50371, 17.5532, 17.95833, 18.39117, 18.33504,
    17.8704, 17.9205, 18.5695, 22.67487, 23.5924, 20.72069, 23.62688,
    19.86155, 18.52993,
  17.45345, 17.47861, 17.45648, 17.50938, 17.48845, 17.46891, 17.47478,
    17.53331, 17.62432, 17.689, 17.78954, 18.16795, 18.43784, 18.8099,
    18.87566, 18.15181, 18.04856, 18.3693, 18.43196, 18.61376, 19.32446,
    20.51937, 21.50186, 21.04949, 25.80162, 28.57952, 23.03765, 23.74278,
    19.86379, 19.02155,
  17.47966, 17.50602, 17.68349, 17.83652, 18.07771, 18.53994, 18.61656,
    18.34947, 18.38627, 18.71038, 18.80992, 19.01122, 18.80091, 18.46768,
    19.28775, 20.15841, 19.59123, 18.66876, 18.87869, 19.21922, 21.40819,
    22.70303, 21.795, 26.18243, 28.15458, 24.58984, 25.42794, 23.28273,
    19.76936, 18.28512,
  17.98206, 17.82283, 18.0812, 18.41018, 18.72165, 18.88528, 18.83246,
    18.69647, 19.21811, 19.62283, 19.38612, 19.23476, 19.07873, 19.32885,
    19.95304, 20.44557, 19.74273, 19.12056, 19.52479, 23.68945, 25.25931,
    20.95239, 20.77768, 22.59639, 24.26248, 23.92978, 23.05892, 23.62772,
    24.12274, 19.95362,
  18.31161, 18.47304, 19.15732, 20.08542, 20.03667, 19.53495, 19.53091,
    19.3834, 19.07294, 19.14297, 19.20079, 20.7396, 22.66089, 22.91166,
    22.36777, 28.90218, 35.60828, 27.78237, 22.3521, 24.0846, 22.67473,
    19.70906, 20.10061, 20.75568, 23.06287, 22.73056, 25.45693, 37.63597,
    33.9181, 19.32213,
  19.12654, 19.49366, 20.20997, 21.06671, 21.16929, 20.9153, 21.68042,
    23.10293, 23.27794, 23.13784, 23.71969, 23.35059, 22.41071, 22.62753,
    27.74721, 34.89346, 32.12399, 24.62015, 22.13958, 21.79696, 20.4387,
    19.61156, 19.99481, 21.94396, 23.36197, 20.96922, 30.05474, 45.16702,
    33.4827, 17.91279,
  20.37374, 20.83632, 21.74624, 22.69891, 22.72483, 24.75036, 26.86819,
    24.86809, 23.29079, 23.16495, 22.89514, 21.94906, 21.04045, 21.21879,
    23.29539, 24.95357, 23.77133, 22.26496, 20.70431, 20.39393, 19.78681,
    19.46564, 20.63316, 22.90666, 22.71892, 21.11987, 32.84111, 38.46326,
    23.70991, 18.11383,
  23.30566, 23.67711, 24.75444, 25.14695, 25.53268, 27.34895, 26.47853,
    24.62427, 24.25084, 23.81627, 22.82195, 21.69011, 21.02002, 24.02868,
    25.78262, 22.54383, 22.38125, 23.98615, 24.20699, 21.82073, 19.75072,
    21.01941, 24.87456, 25.80146, 22.66596, 23.00568, 28.93903, 27.75877,
    20.0158, 18.19356,
  27.34121, 29.22011, 30.72876, 31.98626, 32.01125, 29.04693, 25.21054,
    24.76595, 23.81502, 22.78443, 23.25091, 26.07911, 27.11636, 26.56226,
    25.27828, 25.23518, 26.01204, 26.65122, 25.3393, 23.52651, 23.50718,
    24.10754, 25.09259, 23.73251, 28.45745, 37.46317, 31.09157, 20.77319,
    18.57431, 17.4731,
  40.16173, 43.50003, 39.7831, 34.7798, 33.32797, 31.88383, 28.33571,
    29.71086, 30.71313, 37.24941, 40.87343, 27.68148, 23.82526, 23.24951,
    22.79198, 23.68247, 24.81637, 24.76586, 23.65933, 23.32749, 25.61911,
    25.37193, 22.58071, 20.69561, 24.4453, 28.35162, 23.08371, 18.06163,
    17.74262, 17.30218,
  54.66466, 43.81795, 46.06425, 47.07719, 45.69779, 39.11295, 41.70016,
    38.68387, 31.63508, 35.48743, 34.89762, 22.51383, 23.44475, 24.24513,
    22.47627, 22.88375, 22.34451, 22.19824, 21.87439, 22.4078, 25.1425,
    24.17715, 20.24933, 23.5476, 25.49542, 19.98743, 17.70306, 18.03517,
    17.95215, 17.47323,
  62.07199, 57.46777, 73.91909, 76.6167, 79.16524, 71.3382, 53.99493,
    34.62419, 32.83178, 30.61568, 27.62742, 21.36876, 25.89527, 28.1315,
    23.72847, 22.75569, 22.83967, 22.18084, 21.62796, 23.81321, 25.4657,
    22.53751, 19.88637, 24.70135, 26.12883, 19.2522, 17.90365, 18.19195,
    18.44065, 17.74867,
  66.75662, 76.76749, 78.46954, 78.75067, 72.89565, 63.54493, 58.28893,
    51.76908, 43.10969, 38.2153, 44.13007, 42.93855, 44.98223, 44.11743,
    37.69113, 29.07627, 23.37571, 24.81381, 26.13867, 27.13711, 24.71502,
    23.66298, 25.25241, 22.3794, 20.06834, 18.44925, 17.92208, 17.77752,
    18.15506, 17.71184,
  49.61759, 56.07655, 53.14254, 50.12214, 44.22936, 49.3099, 68.49505,
    65.82857, 56.53954, 56.86963, 55.15599, 42.14478, 32.54387, 37.37976,
    39.06562, 27.13691, 26.55802, 26.60127, 29.29871, 30.51375, 27.1956,
    24.39468, 21.77984, 19.3255, 18.12809, 18.44084, 17.96628, 17.66627,
    17.6862, 17.4582,
  38.83432, 38.14384, 37.27424, 35.77081, 35.25331, 39.8949, 46.3826,
    44.46638, 41.50978, 40.25724, 37.18236, 29.37162, 24.98923, 28.71128,
    28.51245, 26.02494, 27.38538, 25.86999, 26.72003, 26.66781, 22.56797,
    20.41101, 18.52353, 18.4245, 18.64592, 18.42173, 18.04086, 17.78115,
    17.64815, 17.39973,
  35.93325, 34.45142, 33.07785, 32.61, 33.33764, 34.17141, 34.61691,
    34.37091, 33.05849, 30.74479, 26.43608, 25.79642, 29.1024, 27.66783,
    26.35744, 26.24187, 25.68312, 23.9773, 25.12553, 24.16664, 19.08863,
    19.1561, 18.94824, 18.66598, 18.48873, 18.4389, 18.00233, 17.58327,
    17.54907, 17.38856,
  32.29085, 31.55659, 30.89895, 31.35312, 31.65242, 32.31908, 32.5793,
    32.02741, 30.72882, 27.36526, 26.26602, 28.8232, 29.25144, 28.8988,
    30.25105, 28.01467, 24.13759, 21.92969, 24.30918, 23.33173, 19.14032,
    19.49661, 19.34135, 18.91374, 18.133, 18.13193, 17.87324, 17.42827,
    17.39665, 17.31563,
  32.13688, 32.18661, 30.90339, 30.31548, 30.38916, 30.22685, 30.00719,
    29.40564, 27.71345, 25.83239, 27.58306, 27.93654, 24.42842, 25.17608,
    26.02223, 24.85715, 24.36315, 24.64721, 26.72563, 25.72401, 21.84966,
    20.34642, 19.58613, 19.01841, 18.037, 17.85818, 17.72437, 17.42009,
    17.35739, 17.29505,
  32.65219, 32.68618, 30.93769, 29.33722, 29.14268, 28.80381, 28.45414,
    27.85718, 26.82214, 27.78617, 28.31402, 24.52538, 22.17528, 22.21601,
    21.9702, 21.36179, 22.55122, 24.42441, 26.06936, 26.52053, 24.68601,
    22.0129, 19.8211, 19.13098, 18.37928, 17.90452, 17.707, 17.45602,
    17.34257, 17.29314,
  32.19168, 32.02583, 30.21425, 28.66102, 28.24263, 28.13919, 27.99826,
    27.57648, 27.34139, 28.41056, 26.16245, 21.62716, 21.47717, 21.59197,
    21.09291, 20.45091, 20.79756, 21.56184, 22.65369, 23.19153, 23.23401,
    22.93659, 21.44734, 19.74526, 18.73266, 18.14666, 17.69665, 17.45699,
    17.36105, 17.2939,
  32.51933, 31.22673, 29.64949, 28.59502, 28.30639, 27.92588, 27.92945,
    27.4884, 27.85193, 27.4368, 23.39667, 20.38734, 20.72141, 20.82921,
    20.56922, 20.3713, 20.14343, 20.09443, 20.38798, 20.35642, 21.54693,
    21.96307, 21.43983, 21.84543, 20.4889, 18.62468, 17.80397, 17.55672,
    17.37931, 17.30153,
  32.00123, 31.07568, 29.29679, 28.33035, 28.87014, 29.26397, 28.9517,
    27.78994, 27.56469, 25.57249, 21.47713, 20.07298, 20.24083, 20.3644,
    20.10963, 20.46605, 20.42224, 19.60763, 19.30629, 19.30245, 20.50345,
    20.53458, 19.68251, 21.32477, 21.73345, 19.52884, 18.0933, 17.97084,
    17.61176, 17.32605,
  31.48271, 30.78596, 29.96568, 29.6108, 29.76874, 29.90248, 30.23644,
    29.73097, 29.221, 25.408, 21.1344, 20.68292, 20.94173, 21.3214, 21.16815,
    21.1516, 21.22143, 20.38795, 19.42848, 19.39387, 19.73176, 19.54927,
    19.21514, 19.61966, 20.82735, 21.06009, 19.53823, 18.32672, 17.94069,
    17.44358,
  31.36336, 32.09675, 29.96651, 29.24212, 29.58327, 29.52027, 29.22317,
    29.13418, 29.74892, 26.02302, 21.35195, 21.0432, 21.30546, 21.56312,
    21.58048, 21.60597, 21.28165, 20.92842, 20.08161, 19.28812, 19.45027,
    19.55687, 19.4393, 18.97743, 18.92325, 20.22389, 20.30765, 19.04979,
    18.77361, 17.82884,
  31.84781, 33.88553, 32.35243, 30.52207, 29.50103, 28.75316, 29.64378,
    30.61927, 29.09116, 25.12675, 21.95438, 21.48849, 21.74239, 21.50676,
    21.05442, 21.06164, 20.81964, 20.8257, 20.4354, 19.52738, 19.80082,
    19.94304, 19.15166, 18.582, 18.53214, 19.14614, 20.49201, 19.78365,
    18.82548, 17.80417,
  32.75594, 34.49077, 31.79541, 29.79263, 28.97542, 28.36438, 29.86811,
    30.47551, 27.249, 23.72443, 22.18931, 21.72447, 21.59514, 21.28649,
    20.98172, 20.7199, 20.47377, 20.63846, 20.29072, 19.45872, 19.91504,
    21.03672, 21.02669, 20.17383, 19.93616, 20.10206, 22.01047, 21.68972,
    18.81088, 17.34818,
  32.17481, 32.45567, 30.42584, 29.66182, 30.02474, 29.76955, 30.42784,
    29.05645, 25.21623, 23.12057, 21.87826, 21.43068, 21.29709, 21.23946,
    21.54369, 21.22114, 20.46806, 20.41604, 20.74681, 20.86072, 21.5553,
    21.76851, 21.12513, 20.41041, 20.424, 20.56504, 21.12158, 22.95731,
    21.28985, 17.94948,
  29.66946, 28.90263, 29.3559, 30.59892, 31.62246, 32.63412, 31.572,
    27.85625, 24.60889, 22.99834, 21.09174, 20.08599, 19.99785, 20.49025,
    21.32215, 21.56412, 21.50641, 21.89279, 21.47936, 20.69667, 20.69955,
    20.33534, 19.48178, 19.06371, 19.33339, 19.85147, 20.00098, 20.11783,
    20.6685, 18.5001,
  28.59318, 28.72296, 29.02035, 29.11875, 29.531, 31.94436, 32.45645,
    27.91001, 24.26975, 23.16375, 22.16406, 21.75408, 21.78732, 22.23742,
    22.63919, 22.70653, 21.87974, 20.81978, 20.25599, 19.44098, 18.92022,
    18.7878, 18.58056, 18.50018, 18.59423, 19.14065, 19.34761, 18.75641,
    18.28341, 17.53936,
  11.96444, 11.99205, 12.01943, 12.03103, 12.02609, 12.02356, 12.02962,
    12.044, 12.0894, 12.12499, 12.87956, 12.86131, 12.1227, 12.27005,
    12.35559, 12.12531, 12.06655, 12.07981, 12.07665, 12.56379, 12.74235,
    12.32375, 12.27999, 12.66514, 12.82099, 12.49922, 14.7704, 16.00168,
    13.72616, 12.55299,
  12.23164, 12.22766, 12.11437, 12.28881, 12.17665, 12.07459, 12.11325,
    12.1517, 12.20966, 12.34122, 12.72885, 13.17913, 13.35388, 12.74698,
    12.61048, 12.58892, 12.18051, 12.2102, 12.59093, 13.01297, 12.93377,
    12.39243, 12.37835, 12.91546, 16.50642, 16.64264, 15.70138, 18.2586,
    14.6025, 13.11455,
  12.17231, 12.17263, 12.14128, 12.19771, 12.15847, 12.10632, 12.11403,
    12.17191, 12.26291, 12.30945, 12.37334, 12.75708, 13.00186, 13.34279,
    13.3678, 12.6865, 12.62937, 12.88473, 12.87936, 12.99973, 13.5364,
    14.41721, 15.22296, 14.72052, 19.56684, 21.66012, 17.69273, 17.96491,
    14.49192, 13.52417,
  12.12485, 12.12863, 12.26625, 12.37867, 12.60378, 12.99439, 13.00012,
    12.78194, 12.83827, 13.08265, 13.14143, 13.38364, 13.11837, 12.928,
    13.70163, 14.37317, 13.7275, 12.92844, 12.94735, 13.08757, 15.23738,
    16.33972, 15.61203, 19.91488, 21.38368, 19.26395, 20.08937, 17.41082,
    14.29424, 12.94042,
  12.44088, 12.26961, 12.47553, 12.76907, 13.06209, 13.19622, 13.13105,
    12.98555, 13.56753, 13.98792, 13.83184, 13.5517, 13.24837, 13.42355,
    14.02121, 14.34754, 13.41717, 12.86657, 13.15593, 17.39375, 18.53636,
    14.89311, 14.82267, 16.95024, 18.46996, 18.01056, 17.27949, 17.83174,
    18.10794, 14.13062,
  12.45407, 12.51043, 13.17667, 14.08223, 14.06182, 13.54857, 13.47768,
    13.30388, 13.11664, 13.24249, 13.14094, 14.53769, 16.03674, 16.21865,
    15.50498, 21.39781, 26.4648, 19.84945, 15.79244, 18.00773, 16.57281,
    13.76064, 14.24876, 14.80347, 17.29272, 16.71244, 19.16267, 29.38397,
    25.67542, 13.68932,
  12.58986, 12.86694, 13.64742, 14.54253, 14.67614, 14.24563, 14.77742,
    16.13215, 16.28335, 16.2048, 16.86776, 16.47639, 15.67, 15.69851,
    20.24622, 26.76173, 24.78133, 17.97487, 15.91057, 15.71036, 14.44716,
    13.71279, 14.10784, 16.01142, 17.39437, 15.17078, 23.86723, 36.54046,
    25.77203, 12.52189,
  12.83387, 13.16132, 14.03394, 14.83048, 14.77708, 16.77974, 18.62104,
    16.84708, 15.72247, 15.87451, 16.00731, 15.10048, 14.25383, 14.37572,
    16.88127, 18.68281, 17.38977, 15.79061, 14.63014, 14.43318, 13.92824,
    13.66666, 14.65954, 16.76509, 16.62704, 14.78323, 26.72138, 31.06232,
    17.62219, 12.66605,
  14.3983, 14.48275, 15.53292, 15.72087, 16.22342, 18.254, 17.5514, 15.78724,
    15.79881, 15.94233, 15.45602, 14.65669, 14.19039, 17.22344, 18.61804,
    15.94415, 16.10122, 17.38114, 17.27683, 15.28529, 13.68763, 14.69719,
    18.03157, 18.80301, 16.35511, 16.17234, 22.25553, 21.08136, 14.21008,
    12.74155,
  16.81028, 17.94836, 19.59745, 20.80602, 21.15767, 18.59422, 15.58787,
    15.28667, 15.01935, 14.39885, 15.4782, 18.39092, 19.55977, 19.36428,
    18.46599, 18.32403, 18.97055, 19.64144, 18.72472, 17.40176, 17.20446,
    17.97748, 19.13187, 17.81134, 22.20625, 29.88274, 23.94389, 15.1991,
    13.21031, 12.19092,
  26.90789, 29.78289, 27.12157, 22.85136, 22.02756, 21.12844, 18.46453,
    19.89983, 21.12754, 27.71633, 30.04562, 19.80444, 17.29189, 16.84176,
    16.3446, 17.32817, 18.52493, 18.65974, 17.74706, 17.70424, 19.83989,
    19.69753, 17.14855, 15.29353, 19.30796, 23.48061, 18.02516, 12.90424,
    12.42513, 12.0355,
  40.18684, 31.06059, 32.5969, 33.30154, 31.84444, 27.59807, 30.44906,
    28.13438, 22.97673, 27.60127, 26.7968, 15.93684, 16.78069, 17.61878,
    16.53251, 16.9243, 16.562, 16.57768, 16.36837, 17.02039, 19.79797,
    18.69445, 14.87957, 18.1469, 19.86558, 14.73796, 12.4719, 12.71927,
    12.61999, 12.17853,
  45.11911, 41.597, 59.02739, 64.11071, 64.67487, 57.8405, 43.35157,
    26.34664, 24.77231, 23.40252, 20.13347, 14.57025, 19.09548, 21.21033,
    17.64095, 16.99231, 17.10514, 16.56733, 16.15182, 18.55187, 20.21209,
    17.21836, 14.48928, 19.83541, 21.0692, 14.01822, 12.59095, 12.89156,
    13.10168, 12.42342,
  53.46383, 77.33868, 78.53797, 75.29031, 66.6295, 57.00908, 47.61406,
    41.50006, 33.89538, 28.77871, 33.66117, 32.78987, 36.08124, 35.65901,
    30.03837, 22.26621, 17.64394, 19.00683, 20.38784, 21.60154, 19.28032,
    18.37575, 19.83855, 17.43167, 15.07959, 13.15929, 12.64645, 12.52455,
    12.90512, 12.41756,
  39.67617, 47.92122, 46.53112, 44.6105, 38.86863, 41.16177, 55.23615,
    53.84952, 44.63372, 44.72825, 44.66701, 34.03912, 26.03676, 30.84641,
    32.16315, 21.09458, 20.44167, 20.49878, 22.49693, 23.87366, 21.74616,
    19.23761, 17.00697, 14.25593, 12.76327, 13.12838, 12.70145, 12.40105,
    12.43919, 12.19495,
  28.86692, 28.92145, 28.77402, 27.73425, 26.85728, 31.3746, 38.16825,
    36.13888, 33.28241, 33.11867, 30.34357, 23.13442, 18.65918, 22.65381,
    22.63488, 19.97972, 21.44196, 19.81347, 20.25098, 20.44921, 17.55379,
    15.41489, 13.3703, 13.25833, 13.3595, 13.09562, 12.76066, 12.50267,
    12.38798, 12.13418,
  26.79174, 26.00299, 24.83778, 24.13538, 24.62465, 25.63981, 26.30434,
    26.10472, 25.43276, 23.99056, 20.17646, 19.87137, 22.38253, 20.9758,
    20.31205, 20.27608, 19.92254, 18.04823, 18.85603, 17.95475, 13.77423,
    13.8419, 13.69405, 13.47892, 13.248, 13.11837, 12.70512, 12.32607,
    12.30695, 12.12749,
  23.92139, 23.19756, 22.36243, 22.66834, 23.11949, 23.96511, 24.60234,
    24.6746, 23.85234, 21.17225, 20.03629, 22.53433, 23.29769, 22.63993,
    23.97499, 22.09005, 18.41595, 16.23885, 18.38643, 17.28268, 13.72638,
    13.98974, 13.90566, 13.55429, 12.85554, 12.83243, 12.56567, 12.16114,
    12.14864, 12.06339,
  23.51978, 23.44691, 22.27876, 21.97335, 22.35632, 22.64368, 22.9152,
    22.74995, 21.42834, 19.81038, 21.40286, 21.94016, 19.16727, 19.83831,
    20.62506, 19.43524, 18.53406, 18.55049, 20.17015, 18.90111, 15.98022,
    14.75399, 14.01888, 13.55046, 12.68714, 12.5503, 12.43409, 12.14994,
    12.10131, 12.03819,
  23.99884, 24.17653, 22.75395, 21.6013, 21.77927, 21.71252, 21.61227,
    21.31319, 20.50431, 21.52752, 22.19596, 19.0035, 16.90736, 16.91241,
    16.64017, 16.10414, 17.04596, 18.68574, 19.68391, 19.77069, 18.6704,
    16.31951, 14.14511, 13.6195, 13.00409, 12.57923, 12.41338, 12.18832,
    12.10029, 12.03843,
  23.83169, 24.08788, 22.66637, 21.47623, 21.27477, 21.21878, 21.14405,
    20.97651, 20.99743, 22.44226, 20.69789, 16.58176, 16.36251, 16.2114,
    15.56101, 15.00697, 15.32879, 16.09856, 16.74377, 17.01461, 17.58861,
    17.36767, 15.66212, 14.24009, 13.41124, 12.81359, 12.41461, 12.17923,
    12.09443, 12.04078,
  24.49911, 23.82944, 22.49395, 21.66013, 21.34443, 20.95715, 21.12051,
    21.04995, 21.7423, 21.91772, 18.47242, 15.36246, 15.44967, 15.35695,
    15.02337, 14.84631, 14.67267, 14.64127, 14.8829, 14.90802, 16.22755,
    16.37543, 15.60872, 15.89957, 14.76889, 13.14787, 12.46649, 12.25957,
    12.11464, 12.04223,
  24.51604, 23.93488, 22.24649, 21.40296, 21.84683, 22.20592, 22.24088,
    21.51093, 21.71154, 20.37952, 16.64363, 14.90111, 14.81651, 14.82659,
    14.55819, 14.87571, 14.86286, 14.16669, 13.96592, 14.03033, 15.28261,
    15.01008, 13.97284, 15.55357, 15.91179, 13.89855, 12.7321, 12.65543,
    12.34594, 12.06745,
  24.14316, 23.71441, 22.75875, 22.50562, 22.84853, 23.14412, 23.68245,
    23.44355, 23.04135, 19.7765, 16.05536, 15.31927, 15.36424, 15.62803,
    15.44819, 15.52364, 15.58202, 14.76219, 14.02395, 14.1111, 14.36615,
    14.02509, 13.62852, 14.04703, 15.11158, 15.3251, 13.99959, 12.95332,
    12.62626, 12.15697,
  24.20887, 24.78621, 22.89937, 22.45559, 22.96172, 23.04472, 22.86185,
    22.79388, 23.3612, 20.12226, 16.11888, 15.61793, 15.69783, 15.91562,
    15.98175, 15.94877, 15.55754, 15.20443, 14.56916, 14.05893, 14.01727,
    13.98596, 13.92181, 13.54487, 13.59451, 15.02231, 14.99922, 13.64352,
    13.41978, 12.49214,
  24.65201, 26.70614, 25.17618, 23.54769, 22.95797, 22.36156, 22.97932,
    23.76426, 22.60878, 19.43805, 16.63206, 16.03691, 16.06864, 15.81263,
    15.45585, 15.41536, 15.0987, 15.07329, 14.83564, 14.23459, 14.31542,
    14.36922, 13.73601, 13.28515, 13.27029, 13.97168, 15.31501, 14.40853,
    13.53529, 12.5019,
  25.70898, 27.79968, 25.27179, 23.18302, 22.40729, 21.71269, 23.23391,
    23.94425, 21.19443, 18.3053, 16.98788, 16.29845, 15.94562, 15.62068,
    15.27485, 15.03937, 14.80737, 14.8667, 14.70481, 14.1865, 14.40537,
    15.30303, 15.24429, 14.65799, 14.56401, 14.68984, 16.74208, 16.23717,
    13.45578, 12.09641,
  25.6102, 26.31292, 23.89256, 22.73094, 22.9826, 22.67773, 23.55947,
    22.61655, 19.5341, 17.79457, 16.74559, 15.99922, 15.53553, 15.50391,
    15.75075, 15.43169, 14.76307, 14.65363, 15.16796, 15.58012, 15.87216,
    15.82642, 15.40187, 14.95611, 15.09459, 15.15877, 15.9318, 17.74619,
    15.83615, 12.61566,
  23.37199, 22.4646, 22.59538, 23.76058, 24.55534, 25.12606, 24.50601,
    21.47283, 18.85043, 17.56261, 15.8153, 14.74265, 14.56175, 14.87814,
    15.46494, 15.63778, 15.58502, 15.90871, 15.80069, 15.39568, 15.30051,
    14.87912, 14.11103, 13.78242, 14.06021, 14.55905, 14.72115, 14.93355,
    15.49943, 13.14423,
  22.13339, 22.0753, 22.41172, 22.73144, 23.17064, 24.96998, 25.13775,
    21.3562, 18.38197, 17.46818, 16.47644, 16.09376, 16.32873, 16.46781,
    16.4807, 16.56187, 15.89752, 15.10224, 14.73421, 14.03527, 13.58395,
    13.518, 13.30402, 13.21435, 13.31339, 13.8912, 14.12863, 13.49399,
    13.07297, 12.29657,
  9.120263, 9.13925, 9.170859, 9.181655, 9.179828, 9.172775, 9.178283,
    9.186954, 9.214966, 9.22887, 9.935116, 9.923932, 9.229792, 9.368217,
    9.448371, 9.248065, 9.207582, 9.227704, 9.209998, 9.650956, 9.829584,
    9.449829, 9.406404, 9.740018, 9.809867, 9.475572, 11.57029, 12.76179,
    10.77684, 9.693399,
  9.394567, 9.38293, 9.265995, 9.450251, 9.327814, 9.217011, 9.252104,
    9.275243, 9.325982, 9.438755, 9.862522, 10.27092, 10.33913, 9.792317,
    9.681056, 9.669894, 9.32051, 9.345837, 9.68835, 10.11135, 10.04651,
    9.489573, 9.431941, 9.893044, 13.12667, 13.25816, 12.73272, 15.32966,
    11.77942, 10.30871,
  9.361028, 9.349104, 9.297717, 9.362862, 9.288203, 9.214327, 9.225192,
    9.287506, 9.372293, 9.419847, 9.468145, 9.832932, 10.08977, 10.3407,
    10.34542, 9.756098, 9.744256, 9.999277, 9.974121, 10.0169, 10.43792,
    11.24092, 12.01434, 11.39799, 16.284, 18.67889, 14.7539, 15.1387,
    11.64523, 10.6973,
  9.273421, 9.261703, 9.379002, 9.447789, 9.635265, 9.996705, 10.02324,
    9.818515, 9.820191, 10.03911, 10.12364, 10.35226, 10.0939, 9.968841,
    10.69736, 11.28968, 10.72861, 9.996571, 9.896091, 9.884756, 11.92827,
    13.1127, 12.45199, 16.56647, 18.19433, 16.40836, 17.3054, 14.6021,
    11.47506, 10.15054,
  9.539355, 9.353551, 9.533884, 9.787693, 10.08146, 10.28297, 10.19776,
    9.995981, 10.50746, 11.00631, 10.96184, 10.58695, 10.18934, 10.33785,
    10.96896, 11.25587, 10.22381, 9.64337, 9.879019, 13.80207, 15.01446,
    11.85665, 11.7104, 14.10774, 15.47716, 14.8172, 14.43567, 14.91194,
    15.11074, 11.22744,
  9.522016, 9.511637, 10.10505, 10.97862, 11.08996, 10.62218, 10.46238,
    10.28424, 10.15763, 10.31646, 10.16892, 11.35926, 12.69869, 12.8405,
    11.97982, 17.2276, 21.8201, 15.93312, 12.28535, 14.71834, 13.51758,
    10.78193, 11.27224, 11.70903, 14.156, 13.61211, 15.79205, 26.21273,
    22.92749, 10.82711,
  9.555511, 9.804398, 10.586, 11.44344, 11.66214, 11.17656, 11.5093,
    12.77836, 12.88697, 12.70767, 13.27243, 13.08204, 12.41661, 12.28038,
    16.4643, 23.04735, 21.55977, 14.83449, 12.79487, 12.68088, 11.49037,
    10.79669, 11.1361, 12.93536, 14.39091, 12.0473, 20.74674, 34.34086,
    23.55729, 9.594549,
  9.6897, 9.985185, 10.8171, 11.53712, 11.4285, 13.15703, 14.96597, 13.55323,
    12.53756, 12.61194, 12.75195, 11.82654, 10.89471, 10.94386, 13.75264,
    15.8731, 14.40705, 12.6727, 11.67649, 11.51431, 11.03504, 10.76586,
    11.65571, 13.75186, 13.71688, 11.63475, 24.48997, 29.58986, 15.09728,
    9.72792,
  10.7349, 10.81133, 11.79522, 11.91623, 12.31775, 14.60676, 14.21051,
    12.33556, 12.32299, 12.55603, 12.03124, 11.17381, 10.76656, 13.80789,
    15.31361, 12.8178, 13.01823, 14.21039, 14.07853, 12.27268, 10.70269,
    11.62234, 14.85642, 15.70157, 13.38946, 13.15219, 20.18138, 19.0902,
    11.29489, 9.874834,
  12.39008, 13.35967, 15.02452, 16.25849, 16.73018, 14.56128, 11.78172,
    11.4269, 11.37407, 10.82457, 11.86234, 14.80181, 16.04576, 16.07891,
    15.45725, 15.19427, 15.70734, 16.33225, 15.67141, 14.45912, 14.08385,
    14.96772, 16.29876, 15.0774, 19.12929, 26.86255, 21.53891, 12.67245,
    10.44429, 9.343301,
  20.35229, 23.2318, 21.30106, 17.52251, 17.22638, 16.43432, 13.8773,
    15.43633, 16.5076, 22.80876, 25.46803, 16.68811, 14.50618, 13.92784,
    13.3166, 14.38695, 15.66277, 15.79535, 14.82308, 14.83745, 16.99347,
    16.94249, 14.4253, 12.55474, 16.72509, 21.3115, 15.825, 10.20908,
    9.601441, 9.173144,
  32.58527, 24.52953, 25.34457, 25.54568, 24.2222, 20.89587, 23.95907,
    22.60923, 18.49211, 23.67023, 23.46425, 13.11775, 13.74195, 14.4726,
    13.55844, 14.00517, 13.70547, 13.71887, 13.44157, 14.09492, 17.03037,
    15.95561, 12.0807, 15.29999, 17.17392, 12.12702, 9.675116, 9.908928,
    9.806946, 9.32985,
  39.26484, 33.42875, 45.8933, 51.4846, 52.22634, 47.26056, 35.77319,
    20.98627, 20.11819, 19.6354, 16.74138, 11.57726, 15.89068, 17.70659,
    14.62256, 14.05149, 14.20607, 13.67993, 13.25956, 15.71307, 17.47848,
    14.48211, 11.74468, 17.32473, 18.72287, 11.37703, 9.746158, 10.06735,
    10.30058, 9.600402,
  46.04198, 66.53728, 70.29627, 70.51981, 66.18845, 55.25141, 39.38584,
    34.97029, 27.80151, 23.37422, 28.13114, 27.95173, 31.19178, 31.22046,
    26.33986, 19.17455, 14.69345, 16.16333, 17.63782, 18.93806, 16.62214,
    15.58002, 17.15005, 15.01169, 12.60466, 10.37202, 9.81826, 9.687571,
    10.09469, 9.599909,
  32.72252, 41.50846, 42.51064, 42.9723, 38.14358, 37.47175, 47.84369,
    47.58865, 37.48822, 37.38595, 38.63544, 29.54357, 22.75756, 27.56327,
    28.98104, 18.34233, 17.63279, 17.64812, 19.4742, 20.94928, 18.9345,
    16.50119, 14.56069, 11.65071, 9.888808, 10.29148, 9.864049, 9.539991,
    9.58051, 9.354014,
  22.31127, 22.91224, 23.71719, 23.22893, 21.45277, 25.41232, 32.8712,
    30.50286, 27.60052, 28.37519, 26.64017, 19.77915, 15.59658, 19.74372,
    19.81524, 17.19892, 18.84328, 17.05302, 17.295, 17.68954, 14.96592,
    12.75492, 10.6667, 10.53999, 10.54988, 10.2225, 9.884766, 9.632625,
    9.504563, 9.273438,
  20.96363, 20.62518, 19.74841, 18.81665, 18.82558, 19.82801, 20.64755,
    20.37843, 20.28956, 19.87022, 16.72004, 16.54782, 18.95177, 17.78586,
    17.51379, 17.655, 17.48766, 15.46432, 16.07677, 15.26204, 11.013,
    11.02559, 10.93507, 10.80728, 10.45909, 10.2215, 9.828214, 9.467073,
    9.446176, 9.276322,
  18.60745, 17.95685, 17.01866, 17.13221, 17.5606, 18.39061, 19.14436,
    19.50886, 18.88093, 16.75047, 15.9018, 18.83561, 20.26977, 19.73076,
    21.3243, 19.66775, 16.04813, 13.5243, 15.57537, 14.57704, 10.86006,
    11.08811, 11.09746, 10.82677, 10.06548, 9.97582, 9.726522, 9.305273,
    9.297655, 9.216575,
  18.24256, 18.0398, 16.73499, 16.37692, 16.82956, 17.2379, 17.60582,
    17.52221, 16.35078, 15.16043, 17.20797, 18.5465, 16.54578, 17.32662,
    18.18255, 16.99545, 15.92246, 15.4586, 17.00879, 15.85167, 12.9106,
    11.75805, 11.13402, 10.7364, 9.853744, 9.67961, 9.582242, 9.297517,
    9.241783, 9.180388,
  18.61911, 18.58308, 17.1552, 16.08408, 16.28318, 16.22087, 16.13762,
    15.90657, 15.34694, 16.82741, 18.26825, 15.9981, 14.24788, 14.29681,
    14.0072, 13.50183, 14.37231, 15.68684, 16.53917, 16.75526, 15.69288,
    13.35159, 11.24633, 10.79492, 10.13643, 9.691713, 9.55085, 9.32814,
    9.235478, 9.184644,
  18.25237, 18.38489, 17.04926, 15.9417, 15.76748, 15.67072, 15.54514,
    15.49872, 15.96209, 18.09966, 17.24359, 13.79987, 13.74676, 13.51836,
    12.73659, 12.19193, 12.52806, 13.1868, 13.84757, 14.24116, 14.93376,
    14.51618, 12.53707, 11.30423, 10.56018, 9.960185, 9.550762, 9.320582,
    9.238726, 9.184404,
  18.80724, 18.09149, 16.82002, 16.04269, 15.76727, 15.36495, 15.55202,
    15.77587, 17.00736, 18.03896, 15.36376, 12.54865, 12.75864, 12.57903,
    12.12423, 11.92894, 11.80785, 11.83868, 12.14871, 12.13959, 13.50083,
    13.60965, 12.64891, 12.86076, 11.77732, 10.27751, 9.605246, 9.396685,
    9.257389, 9.186296,
  18.88963, 18.15667, 16.56105, 15.76854, 16.21914, 16.62838, 16.85689,
    16.50714, 17.26283, 16.73555, 13.57787, 11.98625, 11.99051, 11.94421,
    11.63991, 11.95417, 11.98346, 11.37951, 11.21799, 11.27306, 12.54025,
    12.19925, 11.09954, 12.64416, 12.9293, 10.98805, 9.875124, 9.798378,
    9.494386, 9.215111,
  18.51938, 18.01731, 17.02385, 16.85323, 17.4016, 17.86935, 18.66626,
    18.79046, 18.71518, 15.94304, 12.76745, 12.26493, 12.34634, 12.5985,
    12.37504, 12.47358, 12.65428, 11.89853, 11.20901, 11.35894, 11.61959,
    11.18519, 10.71064, 11.12454, 12.17448, 12.41823, 11.14214, 10.14529,
    9.805543, 9.307449,
  18.45648, 18.70176, 17.25712, 17.07737, 17.93581, 18.34809, 18.30914,
    18.35997, 18.9997, 16.12651, 12.66522, 12.51869, 12.70419, 12.89113,
    12.92592, 12.9301, 12.63878, 12.31694, 11.73725, 11.32156, 11.2024,
    11.09164, 11.05988, 10.65842, 10.7453, 12.25747, 12.26556, 10.87544,
    10.62784, 9.666491,
  18.76939, 20.36316, 19.45168, 18.3228, 18.14014, 17.95909, 18.50239,
    19.1288, 18.06677, 15.38888, 13.08605, 12.9231, 13.11055, 12.82281,
    12.46382, 12.47506, 12.1605, 12.16842, 12.04349, 11.45402, 11.45147,
    11.51718, 10.9104, 10.43039, 10.39137, 11.1788, 12.59045, 11.61569,
    10.74822, 9.701363,
  19.99876, 21.88894, 20.09275, 18.44202, 17.69503, 17.11588, 18.77345,
    19.32386, 16.49713, 14.17139, 13.50478, 13.26827, 13.05908, 12.65718,
    12.23233, 12.04648, 11.86636, 11.99648, 11.91581, 11.37201, 11.49519,
    12.39073, 12.34497, 11.76216, 11.69515, 11.90652, 13.99252, 13.44085,
    10.64708, 9.276839,
  20.68586, 21.4528, 18.94234, 17.86221, 17.91692, 17.57513, 18.50673,
    17.61833, 14.7465, 13.66824, 13.31028, 12.96468, 12.58296, 12.49376,
    12.67381, 12.38635, 11.81994, 11.77086, 12.31468, 12.72606, 12.97266,
    12.94209, 12.54305, 12.12198, 12.28724, 12.39497, 13.22337, 14.99335,
    13.05347, 9.795359,
  19.04429, 17.99315, 17.8802, 19.08955, 19.43397, 19.50387, 18.97612,
    16.27404, 14.15866, 13.55872, 12.45408, 11.73459, 11.58077, 11.85184,
    12.43686, 12.60006, 12.5851, 12.99429, 13.00375, 12.67988, 12.5701,
    12.08453, 11.27649, 10.94348, 11.24663, 11.74996, 11.92664, 12.302,
    12.84134, 10.34917,
  17.85875, 17.44408, 17.68063, 18.14637, 18.34325, 19.72916, 19.70052,
    16.25165, 13.8991, 13.5458, 12.95185, 12.78815, 13.11386, 13.27547,
    13.32644, 13.46853, 12.94659, 12.30485, 11.97556, 11.2821, 10.8169,
    10.73369, 10.47602, 10.35143, 10.46358, 11.05513, 11.33053, 10.74004,
    10.33039, 9.488754,
  7.973186, 7.990242, 8.027737, 8.04376, 8.041159, 8.032913, 8.033946,
    8.048784, 8.074722, 8.073693, 8.826356, 8.804604, 8.075763, 8.228913,
    8.301059, 8.099843, 8.065825, 8.073874, 8.050611, 8.49502, 8.685183,
    8.311632, 8.268593, 8.605617, 8.617495, 8.245568, 10.42375, 11.6039,
    9.692305, 8.580989,
  8.240397, 8.224304, 8.138191, 8.346025, 8.21322, 8.086993, 8.114165,
    8.136243, 8.190772, 8.297774, 8.866871, 9.263017, 9.222319, 8.695868,
    8.571443, 8.529737, 8.16875, 8.186211, 8.554447, 9.053319, 8.99999,
    8.360863, 8.264357, 8.72563, 11.8404, 11.86042, 12.03428, 14.85131,
    10.98717, 9.291805,
  8.254949, 8.243596, 8.190176, 8.275659, 8.167935, 8.065071, 8.067138,
    8.144966, 8.251398, 8.301143, 8.336456, 8.760351, 9.090086, 9.295654,
    9.274102, 8.622499, 8.559131, 8.829988, 8.873094, 8.932339, 9.260068,
    9.99421, 10.72513, 9.948231, 15.2435, 17.88038, 14.02124, 14.56568,
    10.82322, 9.762511,
  8.14542, 8.132614, 8.253652, 8.308706, 8.476378, 8.862654, 8.924688,
    8.708917, 8.693224, 8.90357, 8.9844, 9.251497, 8.957376, 8.881643,
    9.618178, 10.1886, 9.661987, 8.881861, 8.698569, 8.565697, 10.66709,
    11.93522, 11.23298, 15.33863, 17.35549, 16.11163, 16.99587, 13.99201,
    10.58859, 9.152332,
  8.427786, 8.214849, 8.384894, 8.633775, 8.967027, 9.222965, 9.137258,
    8.893465, 9.40729, 10.01146, 10.00643, 9.537476, 9.018108, 9.143245,
    9.858903, 10.27757, 9.113475, 8.317585, 8.467416, 12.31664, 13.74369,
    10.73859, 10.49609, 13.36986, 14.91531, 14.27579, 14.05585, 14.2558,
    14.16443, 10.08341,
  8.406523, 8.306298, 8.908498, 9.821161, 9.998323, 9.532512, 9.330395,
    9.151492, 9.105335, 9.324688, 9.099261, 10.16458, 11.45925, 11.65539,
    10.70734, 15.45085, 19.93352, 14.39583, 10.79777, 13.67345, 12.5162,
    9.581956, 10.19202, 10.7047, 13.46293, 12.95248, 14.39357, 24.56836,
    21.98381, 9.811668,
  8.343309, 8.572204, 9.418614, 10.40994, 10.74799, 10.11438, 10.2999,
    11.47754, 11.46968, 11.28975, 11.91244, 11.92764, 11.36996, 11.12718,
    14.90214, 21.56951, 20.79576, 13.9054, 11.6144, 11.62283, 10.39721,
    9.689805, 10.11101, 12.05058, 13.62016, 11.06511, 19.71836, 34.33106,
    23.72426, 8.554447,
  8.464287, 8.773671, 9.708517, 10.53137, 10.43358, 12.05094, 13.71771,
    12.32757, 11.35524, 11.4364, 11.75814, 10.73744, 9.574839, 9.447964,
    12.57855, 15.09081, 13.39158, 11.39925, 10.48498, 10.41542, 10.00087,
    9.735346, 10.63392, 12.86546, 12.7661, 10.45902, 24.38854, 30.37938,
    15.07727, 8.663926,
  9.476638, 9.558084, 10.64645, 10.72834, 11.10243, 13.75265, 13.40282,
    11.17222, 11.09307, 11.38163, 10.8078, 9.775432, 9.183266, 12.37968,
    14.07704, 11.56206, 11.81987, 13.10691, 12.98384, 11.20762, 9.627733,
    10.58523, 14.06302, 14.91197, 12.38242, 12.02522, 20.22446, 19.07663,
    10.42406, 8.83382,
  11.29083, 12.17319, 13.99373, 15.32577, 15.86158, 13.62438, 10.71506,
    10.23623, 10.20784, 9.486408, 10.44019, 13.44637, 14.78166, 15.12413,
    14.65647, 14.16282, 14.66838, 15.41647, 14.8589, 13.54839, 12.99366,
    14.06091, 15.70785, 14.46482, 18.06052, 25.5697, 20.76591, 12.05962,
    9.506387, 8.242508,
  18.09793, 21.57708, 20.48086, 16.66916, 16.49985, 15.46808, 12.66739,
    14.21246, 14.77668, 21.23475, 24.35459, 16.07512, 13.81841, 13.07897,
    12.30961, 13.57413, 15.07902, 15.22919, 14.08476, 13.9687, 16.25145,
    16.33897, 13.66257, 11.69719, 16.29738, 21.48144, 15.53992, 9.238517,
    8.458936, 8.022499,
  31.91241, 24.85983, 23.27155, 23.30274, 21.96945, 18.61567, 21.8888,
    21.00739, 16.93223, 22.87137, 23.20269, 12.21393, 12.53416, 13.43263,
    12.74761, 13.28016, 13.01048, 13.04814, 12.65662, 13.28693, 16.48157,
    15.31657, 11.19944, 14.41906, 16.34848, 11.36721, 8.64184, 8.752133,
    8.679135, 8.18564,
  46.20974, 35.26751, 39.00859, 46.2832, 47.76278, 44.47046, 33.91806,
    19.15776, 18.48264, 18.60064, 15.6099, 10.19368, 14.8243, 17.0852,
    14.03587, 13.45579, 13.55344, 12.88518, 12.40097, 15.069, 17.04644,
    13.74697, 10.74851, 16.90524, 18.29098, 10.41294, 8.578108, 8.960989,
    9.21043, 8.458466,
  48.50631, 62.09426, 62.75305, 66.08949, 62.85188, 53.11489, 37.88665,
    32.51153, 25.81437, 21.81191, 26.51559, 26.44118, 30.03406, 29.58419,
    25.38157, 18.64943, 14.15334, 15.66925, 17.193, 18.66379, 16.11411,
    14.98537, 16.68003, 14.64185, 12.03525, 9.313957, 8.69128, 8.60473,
    9.050714, 8.477404,
  30.75446, 38.32033, 39.85477, 42.01938, 37.73629, 36.17255, 45.96858,
    45.94165, 35.06999, 35.55329, 37.70478, 29.19497, 22.37395, 26.7812,
    28.4586, 18.05725, 17.24356, 17.39123, 19.34566, 20.9202, 18.66226,
    16.20483, 14.43999, 10.98366, 8.843101, 9.268702, 8.801624, 8.445057,
    8.514917, 8.235385,
  18.97913, 19.91894, 21.68044, 21.73852, 19.74668, 23.78875, 31.47469,
    28.64258, 25.7361, 27.41834, 26.30486, 19.49404, 15.1559, 19.68269,
    19.61583, 16.96879, 18.78731, 16.92038, 17.18807, 17.77122, 14.92736,
    12.32158, 9.847272, 9.628448, 9.606446, 9.204911, 8.848419, 8.571327,
    8.427026, 8.149386,
  18.0269, 17.98402, 17.43682, 16.32323, 16.02748, 17.22203, 18.30924,
    17.88971, 18.15104, 18.45124, 15.78183, 15.90296, 18.5393, 17.31842,
    17.15838, 17.52629, 17.58507, 15.30749, 16.00204, 15.10706, 10.33991,
    10.21611, 10.02094, 9.858309, 9.50705, 9.183563, 8.740192, 8.378807,
    8.362255, 8.149321,
  15.80329, 15.23163, 14.25775, 14.28075, 14.68487, 15.50716, 16.40626,
    17.05596, 16.73962, 15.0076, 14.51252, 18.14547, 19.85849, 19.19797,
    21.46365, 19.84115, 15.98546, 13.04923, 15.40424, 14.24031, 10.03149,
    10.22613, 10.20199, 9.880954, 9.042871, 8.941072, 8.639755, 8.180474,
    8.188252, 8.083621,
  15.46134, 15.1435, 13.71675, 13.35656, 13.8365, 14.35953, 14.82774,
    14.94881, 14.09539, 13.1877, 15.92665, 17.81463, 15.87195, 17.11567,
    18.53857, 17.18309, 15.75709, 14.91017, 16.73004, 15.31459, 11.94923,
    10.83374, 10.27192, 9.78486, 8.779239, 8.603849, 8.49747, 8.172828,
    8.118608, 8.044846,
  15.86524, 15.61718, 14.06993, 13.0034, 13.27281, 13.32838, 13.37611,
    13.26999, 12.88501, 14.90724, 17.0936, 15.15648, 13.48912, 13.95658,
    13.88884, 13.35355, 14.36588, 15.5604, 16.27515, 16.29706, 14.83187,
    12.48226, 10.43117, 9.845539, 9.079354, 8.597086, 8.435898, 8.200416,
    8.104886, 8.041804,
  15.34489, 15.33849, 14.0039, 12.91619, 12.85612, 12.86055, 12.76376,
    12.74414, 13.46519, 16.35608, 16.08932, 12.97866, 13.20574, 13.12342,
    12.3271, 11.70865, 12.03946, 12.56074, 13.19118, 13.67472, 14.47309,
    13.95959, 11.67715, 10.36649, 9.557898, 8.877638, 8.450761, 8.187799,
    8.100698, 8.04127,
  15.9081, 15.12934, 13.88972, 13.16301, 12.93362, 12.54953, 12.7165,
    13.05644, 14.72898, 16.39538, 14.18466, 11.7355, 12.2149, 12.05475,
    11.44366, 11.06619, 10.81625, 10.84792, 11.29623, 11.32625, 12.91686,
    13.05563, 11.95172, 12.01807, 10.83571, 9.247141, 8.509642, 8.268072,
    8.117218, 8.042681,
  16.17217, 15.29287, 13.73228, 12.99541, 13.44363, 13.80254, 14.11296,
    13.94739, 15.20697, 15.2584, 12.47738, 11.14057, 11.2862, 11.12825,
    10.67225, 10.98002, 11.01198, 10.4563, 10.28917, 10.28076, 11.71803,
    11.32571, 10.27137, 11.93935, 12.13037, 9.967892, 8.764565, 8.687812,
    8.361191, 8.069862,
  15.92484, 15.30054, 14.23444, 14.02483, 14.63548, 15.21237, 16.22216,
    16.812, 17.12764, 14.54189, 11.52106, 11.27061, 11.43122, 11.62729,
    11.3751, 11.58668, 11.82257, 10.98519, 10.20056, 10.32443, 10.65997,
    10.20321, 9.712987, 10.26061, 11.40422, 11.4455, 10.01324, 9.073944,
    8.734544, 8.17349,
  15.82334, 15.71219, 14.44753, 14.43865, 15.51361, 16.28646, 16.57413,
    16.82232, 17.62222, 14.71861, 11.24932, 11.38686, 11.73697, 12.04097,
    12.15341, 12.15788, 11.85595, 11.45257, 10.77509, 10.38284, 10.24913,
    10.11476, 10.14343, 9.698891, 9.786054, 11.41782, 11.30332, 9.819548,
    9.603706, 8.539357,
  15.94274, 16.95111, 16.4422, 15.89472, 16.07546, 16.32482, 16.96925,
    17.49644, 16.30087, 13.71647, 11.49692, 11.71986, 12.20204, 12.06066,
    11.76336, 11.73297, 11.32307, 11.30961, 11.16784, 10.55828, 10.54248,
    10.61784, 9.978705, 9.435372, 9.352304, 10.2489, 11.70842, 10.57041,
    9.751559, 8.596832,
  17.08307, 18.41238, 17.56613, 16.53499, 15.78612, 15.33219, 17.18948,
    17.68344, 14.40604, 12.24556, 11.96908, 12.21008, 12.27212, 11.89964,
    11.41742, 11.18435, 10.977, 11.08651, 10.97668, 10.41965, 10.59712,
    11.52971, 11.39354, 10.78104, 10.78829, 11.03509, 13.23546, 12.44866,
    9.554426, 8.159719,
  18.33663, 18.86809, 16.62811, 16.0455, 16.04628, 15.6463, 16.6533,
    15.58037, 12.43125, 11.72443, 11.95473, 12.07481, 11.82151, 11.66333,
    11.76801, 11.39718, 10.79469, 10.71611, 11.24746, 11.70305, 12.0291,
    12.09361, 11.73572, 11.27577, 11.5036, 11.63791, 12.5748, 14.38398,
    12.14117, 8.667638,
  17.20062, 15.95575, 15.83482, 17.23812, 17.53977, 17.48248, 16.80866,
    13.85388, 11.86029, 11.78169, 11.19201, 10.8063, 10.69058, 10.94342,
    11.55946, 11.61452, 11.51917, 11.94611, 11.99655, 11.77291, 11.75798,
    11.22167, 10.3468, 10.01015, 10.39111, 10.94972, 11.11243, 11.62993,
    12.14217, 9.250672,
  15.91968, 15.40191, 15.87014, 16.34013, 16.42304, 17.73219, 17.44608,
    13.79247, 11.70037, 11.84308, 11.68847, 11.73703, 12.08542, 12.29618,
    12.43559, 12.57452, 12.04892, 11.45662, 11.07029, 10.32365, 9.881734,
    9.779625, 9.466116, 9.337656, 9.495259, 10.16997, 10.45003, 9.730761,
    9.374318, 8.405682,
  8.009446, 8.027488, 8.060293, 8.075423, 8.076065, 8.069081, 8.071639,
    8.088102, 8.097072, 8.084064, 8.746736, 8.820175, 8.096577, 8.240499,
    8.348562, 8.142766, 8.104821, 8.115931, 8.077852, 8.460436, 8.697151,
    8.342929, 8.286453, 8.627042, 8.642935, 8.266115, 10.36364, 11.82166,
    9.853215, 8.759993,
  8.258984, 8.286191, 8.16094, 8.373253, 8.261749, 8.135169, 8.1503,
    8.157874, 8.191864, 8.295834, 8.862666, 9.275068, 9.241674, 8.795953,
    8.597046, 8.595224, 8.211188, 8.205556, 8.545941, 9.069209, 9.070544,
    8.432864, 8.250315, 8.741157, 11.77013, 12.23797, 12.42756, 15.95847,
    11.43042, 9.613825,
  8.295975, 8.300571, 8.218016, 8.326048, 8.219708, 8.091785, 8.08228,
    8.143775, 8.250698, 8.325534, 8.37124, 8.800564, 9.211576, 9.403015,
    9.348823, 8.675032, 8.568644, 8.873458, 8.912688, 9.00372, 9.269643,
    9.942466, 10.6087, 9.980599, 15.13758, 18.70378, 14.83151, 15.96349,
    11.31137, 10.15805,
  8.172634, 8.161917, 8.285286, 8.357689, 8.511924, 8.878792, 8.943918,
    8.725267, 8.682845, 8.866932, 9.00294, 9.322383, 9.094064, 8.972747,
    9.709962, 10.22952, 9.839845, 9.005192, 8.711902, 8.493906, 10.56855,
    12.10255, 11.27653, 15.22921, 17.86654, 16.93958, 18.4632, 15.20314,
    11.0617, 9.448025,
  8.476606, 8.227767, 8.380195, 8.625839, 9.012841, 9.3252, 9.222492,
    8.912312, 9.365931, 10.08826, 10.16816, 9.68539, 9.082846, 9.166603,
    9.974776, 10.49924, 9.330323, 8.264165, 8.319402, 12.09433, 14.19174,
    10.9514, 10.53317, 13.6144, 15.52987, 14.9768, 15.09396, 15.21929,
    15.00749, 10.40586,
  8.445333, 8.279043, 8.832699, 9.754606, 10.11755, 9.739396, 9.40826,
    9.195507, 9.150377, 9.415143, 9.174968, 10.10911, 11.49914, 11.66117,
    10.93138, 14.99446, 19.77772, 14.62837, 10.70834, 13.95282, 13.19421,
    9.61734, 10.27634, 11.02219, 13.87611, 13.71145, 14.46097, 25.31245,
    23.78714, 10.23728,
  8.318702, 8.512605, 9.362628, 10.47749, 10.94847, 10.3346, 10.31046,
    11.59172, 11.61723, 11.30224, 11.83086, 12.07951, 11.61674, 11.22634,
    14.71703, 21.72138, 21.63508, 14.45771, 11.80123, 12.03055, 10.64721,
    9.74081, 10.25825, 12.4138, 14.27753, 11.63002, 19.32819, 35.78008,
    26.50395, 8.827418,
  8.415123, 8.737786, 9.717598, 10.69308, 10.57568, 11.99753, 13.90316,
    12.68292, 11.53918, 11.61707, 12.00015, 11.05938, 9.635938, 9.416434,
    12.61282, 15.74228, 13.93698, 11.68722, 10.66423, 10.567, 10.13403,
    9.852684, 10.84662, 13.38475, 13.39934, 10.76742, 25.06555, 33.85899,
    16.50944, 8.820455,
  9.514121, 9.625193, 10.69125, 10.83053, 11.07765, 14.05047, 13.97411,
    11.3228, 11.13712, 11.52378, 11.00236, 9.775984, 8.96914, 12.15088,
    14.44922, 11.86175, 11.90797, 13.46159, 13.40641, 11.56601, 9.706885,
    10.77598, 14.62426, 15.89504, 12.74011, 12.30188, 21.48371, 21.47635,
    10.65483, 9.008617,
  11.50137, 12.08971, 14.17746, 16.00498, 16.22991, 14.20189, 10.90773,
    10.29401, 10.27913, 9.62134, 10.25884, 13.25677, 14.77106, 15.42788,
    15.1317, 14.4673, 14.98161, 15.97683, 15.5665, 13.99797, 13.24055,
    14.4518, 16.59319, 15.34882, 18.6706, 27.32372, 22.78413, 12.76891,
    9.774669, 8.354087,
  17.42286, 22.4983, 21.88798, 16.89509, 16.65125, 15.87558, 12.8291,
    14.23819, 15.13956, 19.88372, 23.63876, 16.46623, 14.10053, 13.46526,
    12.61815, 14.00498, 15.77308, 16.02094, 14.76953, 14.26591, 16.72101,
    17.06876, 14.40567, 12.04979, 17.1254, 23.48377, 17.27541, 9.580371,
    8.597344, 8.064176,
  33.94986, 27.02713, 23.19904, 21.50622, 20.67627, 16.76575, 21.1489,
    21.65039, 17.08586, 22.43043, 23.53674, 12.46747, 12.68251, 13.72328,
    13.02314, 13.83081, 13.64865, 13.68013, 13.11342, 13.5798, 17.01901,
    16.11253, 11.57047, 14.50515, 17.31897, 12.24126, 8.86488, 8.863265,
    8.785038, 8.250656,
  47.44389, 32.6784, 35.06271, 41.87645, 45.72952, 45.17619, 37.08633,
    19.41623, 19.39105, 19.342, 15.76593, 10.04753, 14.94834, 17.5818,
    14.43876, 13.98252, 14.17949, 13.36892, 12.61132, 15.40414, 17.90025,
    14.25804, 11.01644, 17.219, 19.70441, 10.98184, 8.632299, 9.065137,
    9.358399, 8.595798,
  49.07927, 52.81822, 53.7187, 60.14924, 62.19645, 57.96809, 41.37963,
    33.02505, 27.23821, 21.32432, 25.89314, 26.1739, 31.24212, 30.82942,
    26.51857, 19.64945, 14.68267, 16.31679, 17.79923, 19.71667, 17.25565,
    15.03496, 17.23525, 15.75475, 12.85344, 9.479991, 8.790267, 8.73297,
    9.189363, 8.623151,
  31.05559, 35.6451, 40.08725, 47.85882, 50.13079, 45.1123, 46.6631,
    47.03553, 34.80854, 34.42382, 37.56873, 30.99055, 24.20019, 28.71591,
    30.32096, 19.06485, 18.0255, 18.46789, 20.35437, 22.21406, 19.62341,
    17.04372, 15.51827, 11.84729, 8.892606, 9.342192, 8.897632, 8.554335,
    8.601196, 8.334495,
  19.46449, 22.70084, 27.71862, 30.65744, 28.71077, 27.71585, 32.19731,
    28.96932, 25.30869, 27.904, 27.64233, 21.05898, 15.89054, 21.03083,
    21.01718, 17.68791, 19.81444, 17.96823, 17.87712, 18.87388, 15.98219,
    13.37229, 10.51166, 9.895844, 9.665211, 9.294361, 8.931099, 8.688967,
    8.534512, 8.235085,
  18.29242, 19.53189, 19.94945, 18.41846, 16.44843, 17.05008, 18.42768,
    17.40497, 17.93504, 19.02514, 16.47011, 16.25238, 19.17669, 17.90682,
    17.8667, 18.25604, 18.47492, 16.08827, 16.56118, 16.36302, 11.06842,
    10.632, 10.27126, 10.11528, 9.643691, 9.268846, 8.817471, 8.482159,
    8.456961, 8.228176,
  15.70888, 15.44744, 14.09159, 13.39154, 13.55122, 14.69801, 15.61044,
    16.26301, 16.36013, 14.74785, 14.15473, 18.31247, 20.50368, 19.51438,
    22.71402, 21.09841, 16.90635, 13.59434, 16.08097, 15.41124, 10.34207,
    10.46615, 10.38394, 10.10359, 9.174658, 9.003365, 8.727089, 8.243699,
    8.231735, 8.134969,
  15.15947, 14.71241, 12.84858, 12.32218, 12.83516, 13.34719, 13.87912,
    14.17087, 13.44857, 12.38498, 15.34719, 18.00271, 16.09253, 17.60691,
    20.00077, 18.55492, 16.80791, 15.56808, 17.54197, 16.14039, 12.1149,
    11.04281, 10.41547, 9.937269, 8.881838, 8.670593, 8.577357, 8.224195,
    8.164992, 8.093563,
  15.38439, 14.82957, 13.03642, 11.80611, 12.09861, 12.23003, 12.3863,
    12.32849, 11.8341, 13.89679, 16.78252, 15.21892, 13.56785, 14.46323,
    14.82873, 14.38095, 15.41119, 16.63734, 17.17514, 17.00566, 15.23025,
    12.92566, 10.65462, 10.02071, 9.192815, 8.665465, 8.513837, 8.261429,
    8.159353, 8.098902,
  14.55739, 14.33815, 12.90805, 11.72236, 11.72429, 11.804, 11.67625,
    11.49891, 12.18908, 15.464, 15.98768, 12.95917, 13.5084, 13.718,
    13.03939, 12.4759, 12.83716, 13.34614, 13.80158, 14.32654, 15.08223,
    14.67766, 12.13747, 10.65868, 9.696264, 8.986788, 8.539948, 8.26128,
    8.15808, 8.096145,
  15.06457, 14.03835, 12.78226, 12.03995, 11.87258, 11.39322, 11.40937,
    11.66159, 13.59525, 15.85479, 14.10863, 11.84916, 12.6929, 12.71624,
    12.12114, 11.63029, 11.28788, 11.23159, 11.76268, 11.83979, 13.49853,
    14.02942, 12.45046, 12.43023, 11.08162, 9.428673, 8.60356, 8.346334,
    8.173383, 8.094401,
  15.36908, 14.27921, 12.71384, 11.9103, 12.31803, 12.52325, 12.78843,
    12.68086, 14.39376, 15.11913, 12.46265, 11.38838, 11.80865, 11.72682,
    11.18057, 11.36823, 11.38051, 10.84473, 10.69168, 10.62165, 12.32757,
    12.24197, 10.57829, 12.2853, 12.44217, 10.1661, 8.810742, 8.783719,
    8.432554, 8.118136,
  15.16351, 14.34588, 13.2233, 12.85838, 13.42068, 13.93555, 15.19138,
    16.17786, 16.86092, 14.48742, 11.47379, 11.54317, 11.89841, 12.15837,
    11.82889, 12.01081, 12.30035, 11.44213, 10.55108, 10.65961, 11.23961,
    10.73995, 9.887302, 10.51021, 11.65379, 11.65518, 10.17856, 9.183842,
    8.824373, 8.240442,
  14.97229, 14.70217, 13.31331, 13.18276, 14.35322, 15.39894, 16.0765,
    16.64471, 17.64964, 14.82333, 11.24046, 11.67086, 12.16781, 12.5827,
    12.70576, 12.79115, 12.47408, 11.95912, 11.14625, 10.72312, 10.61892,
    10.37997, 10.37886, 9.94754, 9.977476, 11.63728, 11.55649, 9.963251,
    9.738287, 8.708421,
  14.99918, 15.78978, 15.14889, 14.72022, 15.2653, 15.92664, 16.81835,
    17.5605, 16.33894, 13.77267, 11.43089, 11.94778, 12.67316, 12.70711,
    12.39872, 12.36952, 11.91923, 11.77866, 11.55652, 10.86598, 10.78279,
    10.85864, 10.22134, 9.599171, 9.482242, 10.44142, 11.91857, 10.85134,
    9.959027, 8.825384,
  16.07075, 17.11234, 16.40069, 15.70524, 15.3607, 15.11069, 17.35311,
    18.10453, 14.39597, 11.97689, 11.8544, 12.51267, 12.93953, 12.64997,
    12.02121, 11.67704, 11.44769, 11.5219, 11.40803, 10.74156, 10.83961,
    11.78467, 11.69408, 11.0019, 10.98017, 11.29325, 13.5682, 12.95058,
    9.796373, 8.274159,
  17.48736, 18.01537, 15.71163, 15.54249, 15.83449, 15.52778, 16.74721,
    15.7234, 12.03621, 11.27733, 11.8794, 12.4611, 12.47727, 12.27282,
    12.27335, 11.85315, 11.18531, 11.06762, 11.56555, 12.00865, 12.40728,
    12.56086, 12.2064, 11.67603, 11.80274, 12.01692, 13.04504, 14.8435,
    12.55608, 8.829123,
  16.58221, 15.29397, 15.23543, 17.30885, 17.7683, 17.48706, 16.74514,
    13.48594, 11.14106, 11.35891, 11.21867, 11.12487, 11.10541, 11.32388,
    11.9907, 12.05368, 11.81337, 12.20153, 12.35836, 12.19486, 12.22608,
    11.68237, 10.73214, 10.30909, 10.64769, 11.21465, 11.42869, 12.02986,
    12.56835, 9.578094,
  15.57866, 14.99418, 15.68592, 16.63701, 16.74402, 17.83722, 17.40533,
    13.37679, 11.0016, 11.52569, 11.69352, 11.92419, 12.31399, 12.59377,
    12.84601, 13.00206, 12.42737, 11.79725, 11.4436, 10.63468, 10.12682,
    10.02372, 9.672742, 9.501655, 9.670617, 10.34306, 10.66916, 9.995188,
    9.605547, 8.563463,
  13.45463, 13.49063, 13.51662, 13.53263, 13.52736, 13.52691, 13.52336,
    13.53562, 13.55267, 13.56657, 14.35664, 14.54525, 13.59586, 13.76096,
    13.91641, 13.63749, 13.58288, 13.59387, 13.55598, 13.97939, 14.33066,
    13.93232, 13.85789, 14.26762, 14.30217, 13.86867, 16.11732, 18.36057,
    15.86962, 14.53888,
  13.69391, 13.77998, 13.62311, 13.90212, 13.75985, 13.5775, 13.60443,
    13.60652, 13.65221, 13.83252, 14.47567, 15.02371, 15.02229, 14.48857,
    14.19157, 14.23071, 13.72586, 13.70467, 14.11694, 14.73329, 14.74405,
    14.01298, 13.7557, 14.41413, 17.92173, 19.45832, 18.7229, 23.68222,
    17.77881, 15.62168,
  13.77352, 13.80383, 13.72662, 13.85892, 13.72668, 13.56231, 13.54107,
    13.62098, 13.76777, 13.88729, 13.98978, 14.49102, 14.97005, 15.16315,
    15.15451, 14.35719, 14.12075, 14.55469, 14.60137, 14.70105, 15.02991,
    15.93324, 16.73177, 16.28782, 21.68983, 27.11001, 22.43007, 23.98584,
    17.64626, 16.38827,
  13.67958, 13.67418, 13.82391, 13.93996, 14.14967, 14.63958, 14.68408,
    14.34855, 14.29369, 14.48753, 14.65516, 15.0863, 14.91156, 14.61051,
    15.49773, 16.25144, 15.90758, 14.78409, 14.33509, 14.10236, 16.48296,
    18.58864, 17.57786, 22.30831, 25.91099, 24.44819, 27.5231, 22.95511,
    17.2674, 15.38306,
  14.11697, 13.75947, 13.9719, 14.27102, 14.76975, 15.19179, 15.04862,
    14.63071, 15.16343, 16.20555, 16.40682, 15.6235, 14.7257, 14.96004,
    15.90288, 16.4336, 15.20634, 13.78196, 13.90146, 18.37572, 21.5012,
    17.08021, 16.75723, 20.20339, 22.67718, 22.12299, 22.52099, 23.03537,
    22.64462, 16.59688,
  14.05302, 13.84649, 14.54634, 15.70256, 16.21379, 15.76883, 15.27528,
    15.0341, 14.96565, 15.3176, 15.04669, 16.01383, 17.80054, 17.98015,
    17.42216, 21.67564, 28.01581, 22.37213, 17.09159, 20.76159, 20.08679,
    15.45435, 16.27251, 17.42954, 20.51217, 20.65229, 20.92501, 33.85736,
    33.36496, 16.45021,
  13.86556, 14.13941, 15.21046, 16.62469, 17.31429, 16.59571, 16.29126,
    18.03527, 18.28939, 17.91622, 18.45434, 18.72445, 18.00583, 17.52356,
    21.51801, 29.6268, 29.6546, 21.40162, 18.22477, 18.62007, 16.84093,
    15.57451, 16.28618, 18.96433, 21.21115, 18.47566, 25.68124, 44.80548,
    36.79296, 14.76323,
  13.98165, 14.41796, 15.62546, 16.9158, 16.79728, 18.25891, 20.87082,
    19.69378, 18.06651, 18.21608, 18.58465, 17.47513, 15.56143, 15.36516,
    19.0508, 22.84409, 20.51388, 18.10523, 16.76203, 16.66146, 16.07655,
    15.6935, 16.99433, 20.081, 20.22774, 17.59423, 32.22916, 44.07468,
    24.32308, 14.66304,
  15.35789, 15.57406, 16.75094, 16.97936, 17.26562, 21.19326, 21.4763,
    17.86553, 17.64052, 18.08109, 17.40891, 15.77271, 14.75254, 18.52906,
    21.92307, 18.69732, 18.15867, 20.1237, 20.09433, 17.92802, 15.5449,
    16.90583, 21.54634, 23.20853, 19.1895, 19.30712, 29.4199, 30.50967,
    17.01453, 14.81348,
  17.548, 17.99478, 20.84442, 24.17132, 24.0057, 21.38888, 17.19537,
    16.34798, 16.34349, 15.64551, 16.20553, 19.92161, 21.79913, 22.61177,
    22.09863, 21.3176, 22.10641, 23.19769, 22.52843, 20.43818, 19.72978,
    21.29039, 23.64584, 22.33442, 25.4689, 35.81865, 32.19439, 19.78522,
    15.64174, 13.93857,
  24.51068, 31.60236, 32.38892, 24.94681, 24.48001, 23.60676, 20.24184,
    21.66969, 22.87193, 27.01947, 32.28762, 23.96525, 21.16505, 20.37796,
    19.38573, 21.08032, 23.40127, 23.62797, 21.88909, 20.60503, 23.58717,
    24.30597, 21.13629, 18.23459, 23.62537, 30.82668, 24.5611, 15.44776,
    14.27176, 13.55875,
  43.43314, 36.25406, 32.31184, 28.50581, 28.40234, 23.47156, 27.82413,
    28.42326, 24.16813, 29.93877, 31.43797, 18.48571, 18.85067, 20.37367,
    19.82559, 21.05361, 20.86491, 20.85856, 19.84021, 20.08337, 24.16985,
    23.24282, 17.74662, 20.70834, 24.83837, 19.29738, 14.80042, 14.49974,
    14.41073, 13.78312,
  58.1259, 43.65317, 44.8361, 50.1583, 52.59887, 49.98256, 43.80456,
    36.94909, 42.74817, 30.98174, 21.93131, 17.29803, 22.65314, 24.09014,
    22.09736, 20.90609, 21.2852, 20.31351, 19.07593, 22.3682, 25.56385,
    20.86055, 17.04963, 23.86522, 27.73629, 17.12084, 14.25637, 14.72518,
    15.03389, 14.22483,
  64.4272, 53.85577, 55.69033, 61.6499, 66.44554, 67.22955, 58.06619, 56.056,
    46.40421, 29.91713, 32.68203, 34.63809, 40.38139, 41.35337, 36.40394,
    27.22013, 22.00006, 24.08504, 26.14956, 28.75906, 25.51021, 21.4244,
    24.52737, 22.98217, 19.61122, 15.25154, 14.39427, 14.34012, 14.83436,
    14.27019,
  48.2504, 58.15747, 67.0633, 74.93018, 75.02687, 65.86554, 63.52239,
    64.26971, 42.1582, 40.96684, 48.76688, 42.63494, 35.76522, 37.77043,
    40.43272, 27.73787, 26.36859, 27.07645, 29.78706, 31.86383, 27.33356,
    24.32548, 22.82557, 18.43234, 14.63124, 15.11174, 14.52941, 14.16718,
    14.20214, 13.90401,
  34.52397, 44.75367, 52.5329, 52.33617, 45.1073, 44.99583, 48.97241,
    36.43244, 37.22383, 44.84813, 36.20426, 30.64423, 25.3019, 29.24638,
    29.52781, 26.19964, 28.94646, 26.69461, 25.89729, 27.24425, 23.10093,
    20.12286, 16.98566, 15.81159, 15.4204, 15.1154, 14.65733, 14.34531,
    14.13117, 13.78311,
  25.9696, 27.69671, 28.48158, 24.74029, 21.84811, 25.85022, 28.03113,
    23.24681, 28.70907, 31.30405, 21.72029, 21.80474, 26.32122, 25.17372,
    25.74384, 26.53722, 27.4682, 24.25264, 24.05295, 24.95114, 17.79402,
    16.847, 16.17766, 15.93447, 15.42098, 15.07852, 14.56682, 14.13366,
    14.04024, 13.7782,
  19.46068, 19.53928, 17.48663, 16.16495, 16.64706, 18.28113, 19.22599,
    20.45909, 20.58348, 18.22409, 17.5096, 23.06873, 27.20483, 26.46494,
    32.01177, 30.40431, 25.2714, 20.73992, 23.68342, 23.55196, 16.55077,
    16.63128, 16.30857, 16.02207, 14.93896, 14.75912, 14.47084, 13.82676,
    13.79215, 13.66154,
  18.20232, 17.5668, 14.84302, 13.93624, 14.55303, 15.16969, 15.95725,
    16.30548, 15.28047, 13.83871, 17.74123, 22.32095, 21.17329, 24.08025,
    28.70252, 26.99761, 24.75405, 22.95508, 25.72269, 24.04037, 18.72241,
    17.39223, 16.49946, 15.96525, 14.6485, 14.38288, 14.2848, 13.79554,
    13.6985, 13.59659,
  17.74366, 16.66914, 14.28419, 12.66979, 13.09483, 13.33489, 13.55897,
    13.47075, 12.78264, 15.23795, 19.44496, 18.53815, 17.56274, 20.07938,
    21.67116, 21.69675, 23.13613, 24.75632, 25.24268, 24.94449, 22.49491,
    19.81882, 16.88912, 16.07455, 15.00511, 14.38697, 14.17951, 13.84504,
    13.69455, 13.6127,
  16.24575, 15.64871, 13.79038, 12.27417, 12.31056, 12.52594, 12.44367, 12.1,
    12.82608, 16.92643, 18.43791, 15.51196, 17.38827, 18.94566, 19.11174,
    19.17588, 20.05645, 20.86862, 21.04573, 21.67618, 22.75928, 22.39594,
    18.60436, 16.81592, 15.57488, 14.77256, 14.21015, 13.85966, 13.70023,
    13.60882,
  16.82115, 14.98051, 13.49538, 12.50899, 12.43066, 11.91646, 11.90982,
    12.08177, 14.4093, 17.53448, 16.07202, 14.06268, 16.57892, 17.89943,
    18.10853, 18.10145, 17.95776, 17.84905, 18.50579, 18.82497, 20.7249,
    21.55818, 18.98471, 19.0305, 17.38603, 15.41349, 14.31276, 13.97573,
    13.73551, 13.62169,
  17.12531, 15.15188, 13.35284, 12.29499, 12.92721, 13.20045, 13.36874,
    13.10312, 15.2504, 16.64949, 13.95798, 13.59293, 15.60495, 16.84104,
    17.05912, 17.73067, 17.85414, 17.2092, 17.17162, 17.24174, 18.91719,
    19.05081, 16.90778, 19.00366, 19.20364, 16.43729, 14.57788, 14.52888,
    14.05477, 13.64966,
  16.82752, 15.22516, 14.03907, 13.54161, 14.17165, 14.63735, 16.2949,
    17.85006, 18.78653, 15.99357, 12.77169, 13.94035, 15.80462, 17.35967,
    17.85635, 18.48791, 18.90101, 18.00004, 16.97312, 17.16974, 17.88016,
    17.1549, 16.00871, 16.97203, 18.37128, 18.18262, 16.30621, 15.03468,
    14.55406, 13.82202,
  16.33625, 16.1303, 14.25907, 13.74083, 15.17347, 16.64948, 17.78436,
    18.86872, 20.01187, 16.72695, 12.62202, 14.21671, 16.12669, 17.90186,
    18.92681, 19.60599, 19.36631, 18.67718, 17.58648, 17.00869, 16.96879,
    16.60717, 16.6433, 16.263, 16.1586, 18.00595, 17.92838, 15.97703,
    15.6019, 14.44473,
  16.46467, 17.68511, 16.644, 15.86213, 16.52738, 17.6037, 19.01805, 20.2113,
    18.61699, 15.74109, 12.96451, 14.51318, 16.62214, 18.02135, 18.64897,
    19.27482, 18.83397, 18.34327, 17.88926, 16.92074, 16.91885, 17.1683,
    16.44687, 15.54456, 15.31019, 16.5158, 18.14212, 17.03806, 15.81323,
    14.56484,
  17.70328, 19.03544, 18.22662, 16.96834, 16.79642, 16.92496, 20.17372,
    21.49929, 16.54591, 13.50032, 13.46364, 15.04884, 16.85089, 17.91514,
    18.2591, 18.44162, 18.12868, 17.97379, 17.70634, 16.77278, 17.09767,
    18.22603, 17.9614, 16.96927, 16.95712, 17.46498, 19.91532, 19.43092,
    15.64813, 13.83216,
  20.11811, 21.78539, 17.16876, 16.51636, 17.33155, 17.46494, 19.42788,
    18.65981, 13.63334, 12.46107, 13.45202, 14.94841, 16.33767, 17.53398,
    18.55648, 18.55667, 17.70448, 17.43661, 17.82303, 18.15304, 18.95156,
    19.36094, 18.72346, 17.93567, 17.95361, 18.34528, 19.54532, 21.58058,
    19.0575, 14.56959,
  19.00443, 17.39314, 16.69889, 20.52743, 20.84229, 19.69054, 19.29856,
    15.52544, 12.17858, 12.40479, 12.63298, 13.35621, 14.72004, 16.36047,
    18.1246, 18.69519, 18.41006, 18.77784, 18.8323, 18.53271, 18.78321,
    18.23181, 16.97987, 16.3571, 16.73161, 17.43495, 17.7749, 18.62042,
    19.10221, 15.6034,
  17.56341, 16.38657, 18.3643, 21.29276, 20.88394, 20.9387, 20.20131,
    15.34067, 12.05417, 12.74043, 13.27475, 14.38362, 16.1742, 17.83979,
    18.98736, 19.58307, 19.07557, 18.33939, 17.78818, 16.76466, 16.19072,
    15.98214, 15.56112, 15.35343, 15.61266, 16.40986, 16.80555, 16.1083,
    15.58175, 14.27902,
  17.69383, 17.78788, 17.85628, 17.90501, 17.89104, 17.89054, 17.88981,
    17.92297, 17.97192, 18.19475, 19.67476, 20.18002, 18.14319, 18.44797,
    18.76671, 18.13259, 17.9824, 18.05165, 18.06764, 18.72536, 19.37243,
    18.88434, 19.15894, 20.15032, 21.12529, 21.73411, 26.10675, 30.1371,
    23.05617, 19.88801,
  18.29195, 18.55884, 18.1584, 18.69447, 18.39471, 18.02557, 18.1006,
    18.15976, 18.3288, 18.78205, 19.7893, 20.82355, 21.07387, 19.97247,
    19.18596, 19.41889, 18.38052, 18.53541, 19.49366, 20.49478, 20.06165,
    18.93333, 19.65143, 22.98554, 30.34706, 34.19648, 31.16445, 37.88083,
    25.65475, 21.53991,
  18.33304, 18.41099, 18.3002, 18.44939, 18.20907, 18.00248, 18.04214,
    18.22663, 18.48257, 18.66507, 18.96756, 19.83573, 20.55894, 21.09289,
    21.28768, 19.7012, 19.49389, 20.44608, 20.31516, 20.66265, 22.12452,
    25.39083, 28.21387, 30.36439, 39.67225, 46.50235, 38.86309, 38.19417,
    25.52217, 22.86157,
  18.21263, 18.28322, 18.60102, 18.95995, 19.36213, 20.20001, 20.2679,
    19.61917, 19.55692, 20.16939, 20.74196, 21.2298, 20.89339, 20.36002,
    22.44916, 24.20648, 23.23956, 20.64714, 20.24826, 21.39874, 27.10748,
    31.93032, 30.70052, 39.61123, 47.94629, 42.05531, 46.45134, 35.82886,
    24.9579, 20.81603,
  19.11303, 18.47629, 18.99303, 19.64837, 20.59207, 20.97058, 20.61365,
    20.281, 21.60659, 23.31632, 22.88209, 21.62525, 20.73696, 21.71813,
    23.23093, 23.51635, 21.87217, 20.28127, 21.96286, 30.24327, 35.92158,
    28.77472, 29.61063, 34.38667, 36.78274, 36.12222, 35.11362, 37.40295,
    34.8655, 22.3309,
  18.87477, 18.97402, 20.72402, 23.00399, 23.08796, 21.99211, 21.51175,
    20.97797, 20.79083, 20.99586, 21.01847, 23.80928, 28.39999, 29.09592,
    31.73637, 37.57522, 43.26517, 37.13875, 29.46399, 34.16839, 32.18581,
    25.25071, 27.17536, 29.60433, 32.47361, 32.38409, 35.93924, 55.29726,
    48.8585, 21.70741,
  19.05477, 20.20347, 22.61118, 25.02273, 24.70288, 23.0649, 24.54653,
    28.90608, 29.64138, 28.98942, 30.09575, 30.04681, 28.25388, 28.76516,
    35.78043, 46.25546, 43.88876, 35.36523, 29.38565, 29.75628, 26.74705,
    24.51492, 26.39866, 31.673, 36.31139, 37.5195, 47.33755, 61.87315,
    50.59406, 19.62434,
  19.51654, 21.10105, 23.62907, 25.7025, 25.28673, 28.84255, 35.05181,
    32.2197, 28.60928, 29.23576, 28.94909, 26.40096, 23.59039, 25.35213,
    30.54431, 34.97625, 32.60486, 30.19786, 25.84752, 25.53982, 24.41066,
    24.14359, 27.69197, 33.5061, 35.23595, 36.08392, 51.81869, 62.56708,
    37.8899, 19.76963,
  21.93979, 22.6038, 24.82973, 26.31011, 28.67685, 34.17163, 32.2425,
    27.68991, 28.49623, 28.07397, 25.71713, 23.02679, 22.91567, 31.43063,
    38.66624, 31.27057, 29.14505, 31.79852, 31.73892, 28.04962, 23.73458,
    27.77461, 36.97116, 40.25856, 33.04573, 35.82523, 48.61056, 48.73569,
    26.88762, 20.00967,
  26.53127, 32.30302, 35.76888, 38.25237, 40.10259, 35.62941, 23.76096,
    23.38983, 22.62047, 22.36162, 25.36625, 34.61155, 38.92248, 37.88446,
    34.54844, 33.52156, 35.17458, 37.33097, 34.67633, 29.52237, 30.08008,
    32.65084, 36.22237, 37.88622, 46.89619, 60.28094, 52.04884, 29.17663,
    20.87176, 18.35946,
  40.82146, 47.20649, 49.00083, 44.08465, 43.11066, 36.52966, 28.40914,
    32.15144, 36.22277, 43.25626, 51.45668, 37.92965, 32.26307, 30.35168,
    29.18866, 31.73968, 34.74582, 34.65975, 31.91276, 29.40812, 33.46956,
    34.58038, 30.69486, 29.08817, 36.32866, 42.50648, 32.67481, 19.94046,
    18.89644, 17.79334,
  62.16689, 49.93034, 49.35648, 49.54507, 46.82018, 36.83292, 44.7308,
    47.01836, 42.5688, 45.37579, 42.43786, 27.57459, 28.44134, 30.42865,
    30.1325, 32.15325, 31.67131, 30.75749, 29.27023, 30.65994, 34.55484,
    32.42038, 25.34369, 29.78623, 35.52145, 26.44747, 19.44233, 19.19507,
    19.11593, 18.17824,
  76.06164, 63.32627, 75.42687, 83.24338, 84.3484, 78.13108, 65.74779,
    47.63747, 49.28221, 39.12027, 30.38476, 25.9203, 33.74421, 38.57426,
    36.41774, 32.87133, 32.37245, 30.47776, 29.26132, 36.7006, 39.78822,
    28.80123, 25.4125, 32.29221, 36.02269, 22.53422, 18.73514, 19.60183,
    19.88179, 18.80227,
  85.44009, 95.36234, 99.16476, 101.7836, 96.28182, 88.77003, 78.34555,
    70.91833, 55.02068, 42.82193, 53.0102, 55.50667, 61.83736, 63.32521,
    55.44136, 42.19365, 33.80323, 37.05491, 40.81023, 43.9719, 38.40777,
    30.93619, 35.05408, 30.37348, 24.31759, 20.20961, 19.14218, 19.01018,
    19.52582, 18.84058,
  80.77959, 80.49815, 85.47379, 83.50684, 72.8909, 71.66926, 85.25787,
    80.6256, 65.15607, 67.85472, 72.35973, 62.6956, 56.48151, 61.57505,
    59.28043, 44.57879, 42.78306, 45.38028, 50.02755, 50.98537, 41.34271,
    37.75076, 32.38739, 23.7502, 19.57148, 20.07216, 19.31198, 18.76914,
    18.72029, 18.31174,
  73.4229, 73.70982, 73.12894, 66.76898, 66.26524, 73.14329, 80.88202,
    82.46834, 58.69816, 62.58308, 60.88839, 50.07166, 44.04636, 50.90618,
    48.78334, 45.24624, 48.23688, 46.16973, 46.3672, 45.69129, 33.98175,
    28.50587, 23.84414, 21.21237, 20.61972, 20.11102, 19.38297, 18.96344,
    18.61576, 18.14456,
  64.50678, 60.08398, 53.10798, 49.55753, 51.6153, 53.39809, 58.10033,
    63.36027, 48.49874, 48.65784, 43.46096, 41.33825, 46.53109, 42.82455,
    45.95377, 45.82489, 45.65753, 41.43833, 41.98658, 40.39289, 24.9618,
    22.14745, 21.67831, 21.80165, 20.63457, 20.06209, 19.32172, 18.60329,
    18.43956, 18.14132,
  48.65956, 43.43044, 37.70028, 37.46584, 39.82619, 44.26373, 47.31517,
    46.22583, 41.52144, 36.77521, 37.49649, 46.71186, 50.64357, 49.38843,
    54.94143, 49.60199, 40.62672, 35.60634, 40.24137, 36.40557, 22.51321,
    23.20023, 22.9644, 22.11646, 19.81348, 19.54288, 19.1935, 18.18992,
    18.11343, 17.95313,
  39.88219, 36.77192, 31.79497, 31.0056, 35.40847, 39.27235, 37.83455,
    34.77513, 31.29769, 29.78988, 38.80739, 47.52417, 43.4866, 47.1941,
    48.64756, 41.28501, 38.8227, 40.67569, 43.89608, 38.58883, 27.32847,
    26.03606, 23.99742, 21.9416, 19.35518, 19.00581, 18.83215, 18.1257,
    17.99427, 17.87971,
  35.46005, 34.15335, 30.4116, 28.22223, 31.98392, 32.65685, 29.37434,
    26.776, 26.04077, 33.53151, 42.57182, 39.74625, 37.30082, 39.43119,
    36.74973, 33.14037, 34.84164, 40.32352, 42.50137, 41.50496, 35.64764,
    29.98253, 24.54159, 22.03875, 19.95399, 19.05601, 18.68092, 18.23238,
    17.98757, 17.88465,
  33.17589, 32.93055, 28.53673, 26.45215, 28.10458, 27.40684, 24.70824,
    23.93188, 27.49499, 37.01716, 39.27903, 32.58518, 34.83116, 33.67665,
    30.58847, 29.73829, 31.78159, 35.06262, 37.01501, 37.63806, 35.52168,
    32.54398, 27.17114, 22.99963, 20.62733, 19.65256, 18.74953, 18.27279,
    18.0254, 17.89703,
  33.53024, 31.61153, 27.77231, 26.04206, 25.96568, 23.5364, 23.11758,
    24.70262, 31.12625, 37.37486, 33.55468, 29.13336, 31.06282, 29.04861,
    27.48308, 28.24673, 30.225, 31.54836, 32.02912, 31.66243, 31.59102,
    31.09717, 28.11008, 27.09541, 24.13411, 20.92525, 18.9854, 18.50143,
    18.06945, 17.91276,
  32.65051, 31.3563, 26.77516, 24.16697, 25.00356, 25.39868, 26.32809,
    27.1395, 32.41438, 35.12411, 28.45629, 26.07383, 26.65545, 26.16389,
    25.58964, 27.8899, 30.22674, 29.51185, 28.53934, 27.94274, 28.53975,
    28.09488, 25.90069, 27.9706, 27.56162, 22.74931, 19.4968, 19.4295,
    18.61686, 17.97956,
  32.14835, 29.77128, 27.42352, 26.73922, 27.88974, 28.81393, 31.50818,
    32.29894, 35.71831, 33.31701, 25.21289, 24.64174, 25.48357, 26.78081,
    27.88313, 30.26698, 31.8706, 30.20434, 27.96597, 27.12978, 26.47591,
    25.47395, 24.90126, 25.94354, 26.99881, 25.82896, 22.65349, 20.31529,
    19.32597, 18.25997,
  30.1003, 31.33055, 26.84662, 26.5403, 28.9226, 30.57618, 32.21658,
    33.40171, 37.82834, 33.62543, 23.51512, 24.45115, 26.51024, 29.09617,
    31.0488, 32.99321, 32.60144, 30.88762, 27.72129, 25.02049, 25.11847,
    25.53881, 25.14487, 23.74346, 23.06416, 25.10474, 24.78524, 21.76119,
    20.86178, 19.27224,
  31.27805, 34.56981, 30.84181, 29.48611, 30.59143, 31.35526, 33.03069,
    36.08528, 37.10697, 30.48557, 23.65546, 25.43079, 28.61832, 31.02787,
    31.69723, 32.48168, 31.49785, 29.54736, 26.48441, 23.70375, 25.42804,
    26.54107, 23.81426, 21.24763, 20.89608, 22.73764, 24.78525, 23.27742,
    21.13102, 19.49199,
  34.67887, 37.65141, 34.43937, 32.03327, 32.25351, 31.2863, 34.4747,
    36.96997, 33.1594, 26.03934, 24.96186, 27.74401, 30.51762, 31.4921,
    30.98802, 30.59068, 29.4622, 27.76095, 25.31094, 23.28923, 25.35222,
    27.32167, 25.62961, 23.37429, 23.04877, 24.04845, 27.11498, 26.50241,
    20.95811, 18.34358,
  38.39847, 40.41493, 33.73233, 32.55208, 34.87975, 34.45688, 36.16265,
    34.54875, 27.3158, 24.82256, 26.7374, 29.63182, 31.10948, 30.91528,
    30.71933, 29.91345, 27.81321, 26.13762, 25.15396, 25.23575, 28.1937,
    29.39834, 26.83236, 24.89775, 24.43429, 25.36708, 26.84226, 29.1022,
    25.66399, 19.39804,
  34.56688, 30.2878, 30.7167, 35.85878, 38.46073, 39.95967, 37.82608,
    30.08282, 23.9658, 25.63475, 27.13418, 28.01498, 28.3101, 28.35359,
    29.40383, 29.55802, 28.7099, 28.38774, 26.86504, 25.87082, 27.45443,
    26.64371, 23.84542, 22.44377, 22.85695, 24.01657, 24.53894, 25.26859,
    25.27714, 20.8615,
  31.0426, 29.63198, 33.61375, 35.9766, 35.46799, 38.35758, 39.29539,
    29.43039, 23.81232, 26.62209, 28.28194, 29.84976, 30.0518, 30.20247,
    30.94516, 31.35962, 29.96181, 27.42213, 25.1821, 23.32796, 22.71355,
    21.91373, 21.06734, 20.75084, 21.25267, 22.36119, 22.80989, 21.81355,
    20.66122, 18.81504,
  17.39325, 17.70076, 18.10341, 18.50306, 18.60141, 18.92301, 19.36596,
    19.95638, 20.79313, 22.26616, 25.11746, 25.29326, 20.11724, 21.1257,
    21.46991, 20.23488, 20.61009, 21.91075, 23.71399, 26.81769, 28.84387,
    27.56898, 29.26681, 32.97245, 36.13428, 38.0593, 45.30172, 48.78689,
    27.18151, 20.25378,
  20.94196, 21.70935, 20.8721, 22.37758, 21.7403, 21.35088, 22.12965,
    22.80105, 23.78905, 25.0798, 27.03506, 29.27177, 29.97104, 27.03384,
    25.6943, 27.15108, 26.07011, 28.64057, 32.25412, 35.45109, 36.40967,
    37.33287, 40.83728, 49.18869, 57.15123, 53.63327, 47.50715, 51.55973,
    29.02085, 22.64199,
  19.92379, 20.12937, 20.44722, 20.95251, 21.18489, 21.56812, 22.10308,
    22.88925, 23.94639, 25.07942, 26.61245, 29.09816, 31.40755, 34.21114,
    36.65867, 34.93972, 37.54805, 42.02534, 45.34045, 50.96514, 59.26962,
    67.9233, 71.91145, 74.57565, 76.10722, 68.58417, 61.44897, 49.32986,
    29.47507, 24.66115,
  21.82287, 22.8358, 24.78023, 27.01781, 28.98458, 31.42232, 31.8349,
    31.28407, 32.25885, 34.35537, 35.67109, 37.01036, 38.27001, 40.16395,
    47.99741, 53.60808, 52.50491, 51.07724, 57.37523, 65.26818, 76.1105,
    78.63533, 74.44926, 81.77444, 81.48877, 77.5311, 67.72444, 47.5673,
    28.85863, 20.99656,
  27.08212, 26.68488, 29.68081, 31.90467, 33.71545, 33.52235, 33.25255,
    33.83043, 36.46027, 38.7132, 37.85958, 39.25352, 42.34214, 47.94582,
    53.52602, 57.50898, 57.78401, 55.39326, 61.45321, 71.54955, 73.31951,
    61.21114, 61.42359, 70.36028, 76.67738, 74.58709, 65.95274, 69.88464,
    59.0722, 29.78634,
  28.4556, 31.16192, 35.49241, 39.8462, 38.68164, 36.26905, 37.86774,
    39.61263, 41.68371, 47.22481, 55.82129, 69.77067, 84.3538, 84.659,
    88.9883, 94.4514, 93.68252, 83.44162, 70.19693, 69.79153, 62.15596,
    51.86981, 58.69949, 66.30129, 74.36638, 74.50578, 71.11176, 85.30429,
    69.89607, 28.0216,
  32.32626, 37.45927, 43.74879, 50.71568, 54.49327, 59.59483, 70.26276,
    81.69292, 84.8176, 84.99429, 86.09711, 82.32719, 72.82039, 73.47432,
    75.56081, 77.0226, 75.88937, 66.99678, 56.16577, 57.37513, 53.90881,
    53.37802, 59.88037, 69.01552, 71.95474, 63.5471, 67.5341, 77.856,
    57.84277, 19.50761,
  40.12881, 48.37453, 57.00393, 66.17314, 71.27013, 81.84531, 89.52289,
    73.68864, 61.82076, 61.11559, 56.42532, 50.88483, 45.73565, 47.12481,
    49.7923, 54.31961, 56.64714, 55.25684, 48.42236, 49.76581, 49.70551,
    52.7897, 61.12687, 67.94897, 64.20374, 60.95602, 72.16306, 71.05635,
    44.8916, 20.49175,
  55.06586, 60.96079, 67.03669, 70.38974, 70.45184, 73.68254, 62.4964,
    54.21074, 55.52298, 54.53688, 53.04049, 53.01793, 57.21112, 71.27307,
    80.1203, 63.44566, 65.35074, 71.4874, 70.6209, 63.45399, 60.08768,
    74.07495, 88.7198, 88.26905, 72.92682, 80.04671, 80.75103, 63.75866,
    28.88674, 20.33718,
  79.44016, 88.92307, 86.02637, 88.88553, 79.38115, 66.7561, 47.8546,
    56.9795, 60.55367, 71.52502, 84.98264, 99.26937, 96.82527, 91.64101,
    83.68592, 89.94009, 94.0128, 92.43749, 85.33279, 82.1485, 90.53461,
    91.61274, 88.32539, 77.11663, 82.8413, 94.23164, 75.80333, 38.6069,
    20.10715, 16.64207,
  99.62478, 97.83498, 97.27305, 85.61465, 96.76172, 97.65044, 96.25284,
    103.8216, 105.9704, 107.5988, 105.847, 76.84095, 72.36554, 71.52283,
    74.48102, 81.0157, 85.72937, 84.55119, 80.58064, 80.67551, 91.05853,
    85.39552, 64.48431, 55.6471, 62.19512, 60.48209, 37.62776, 20.62914,
    18.93702, 16.34165,
  99.9413, 89.98835, 99.96452, 102.089, 103.8118, 99.04779, 102.1916,
    95.45506, 84.28009, 72.04893, 62.71624, 57.21236, 63.88502, 70.13844,
    72.82289, 73.71999, 72.16561, 70.65137, 66.99392, 67.65341, 75.5659,
    67.49513, 49.08157, 57.5334, 60.08108, 38.96684, 19.48138, 21.58089,
    19.97306, 17.64036,
  106.2439, 107.5143, 111.4743, 112.691, 111.6854, 106.9549, 97.44373,
    84.54823, 85.92252, 63.61077, 62.13036, 65.51649, 77.19632, 86.17336,
    82.72975, 69.8726, 70.19443, 66.56848, 63.2989, 68.94889, 71.30508,
    58.33996, 49.72269, 49.57728, 45.14616, 30.49823, 21.27991, 23.30348,
    22.17396, 19.30879,
  110.7698, 112.1647, 111.1681, 108.5077, 105.1634, 102.101, 100.8459,
    101.0095, 98.4635, 98.69683, 100.7836, 99.97138, 102.8218, 104.2108,
    101.1504, 86.44768, 85.38789, 91.03729, 95.0907, 89.73856, 72.27032,
    53.6056, 48.86682, 35.91015, 28.36945, 25.16933, 21.78897, 20.73967,
    20.52729, 19.03865,
  104.7541, 103.0656, 101.2451, 99.63239, 98.8565, 100.4837, 105.2138,
    106.2627, 103.0344, 103.889, 103.2342, 103.0592, 104.5224, 104.5494,
    102.6766, 101.3673, 100.2534, 101.1608, 100.5306, 87.26443, 54.92908,
    46.5256, 34.02781, 27.7142, 25.22684, 23.86623, 21.18551, 19.49285,
    18.4428, 17.50653,
  100.0192, 100.0632, 100.2043, 100.3754, 101.1356, 104.1315, 107.1524,
    105.3205, 103.5293, 103.3783, 103.4486, 101.6819, 100.9104, 103.2188,
    102.021, 100.9172, 100.8356, 86.60457, 75.38543, 61.52557, 37.85258,
    34.95232, 27.84625, 26.55723, 25.46345, 23.25817, 20.70449, 19.57849,
    18.34701, 17.29216,
  87.42657, 84.96143, 88.69757, 93.40657, 98.07668, 101.9975, 102.8636,
    103.2321, 99.83696, 97.54865, 91.18857, 101.6643, 104.6028, 102.6299,
    101.6061, 93.91188, 81.1692, 67.06478, 61.71397, 54.06252, 31.87735,
    32.88665, 28.52866, 26.54039, 24.48706, 22.94287, 20.27392, 18.27246,
    17.7168, 17.16818,
  70.44382, 74.65971, 75.45348, 79.61593, 82.51398, 86.3611, 88.28549,
    89.06464, 90.4598, 91.03098, 102.6836, 106.6326, 106.3739, 105.2704,
    104.6892, 88.98778, 64.56483, 55.6407, 60.62059, 53.55852, 33.19589,
    33.96243, 29.64048, 27.31628, 22.90043, 21.04584, 19.66361, 17.18,
    17.0001, 16.6556,
  78.31427, 76.52289, 67.53461, 63.82836, 66.6907, 69.07065, 72.89581,
    78.52036, 83.50802, 93.8979, 103.9943, 104.2455, 93.58542, 91.78391,
    84.25964, 74.91439, 74.48502, 77.48172, 78.22774, 64.96249, 42.53582,
    36.13042, 30.46081, 26.39558, 21.46402, 19.51851, 18.64255, 17.1501,
    16.77861, 16.58427,
  75.42455, 69.1373, 58.50254, 51.81567, 55.21263, 59.61218, 66.47066,
    74.40601, 83.66643, 96.98164, 99.89737, 78.22035, 70.1077, 68.29272,
    65.0619, 65.82224, 71.51727, 76.9627, 75.17113, 68.29652, 53.8903,
    42.23124, 31.72342, 26.74676, 22.58359, 19.61554, 18.49052, 17.29665,
    16.71275, 16.5798,
  66.20503, 59.20974, 49.61149, 45.93617, 50.41279, 56.9411, 63.76792,
    70.48021, 77.5891, 83.31723, 73.81082, 56.60619, 62.01212, 62.53341,
    61.90412, 61.65206, 63.39845, 63.05733, 61.15274, 56.77322, 50.63277,
    47.08832, 38.38892, 30.03763, 25.10489, 21.24504, 18.59902, 17.3599,
    16.70647, 16.58194,
  64.55781, 53.13038, 48.02995, 47.0702, 52.25914, 55.13837, 61.495,
    65.09604, 70.85143, 71.39807, 57.73194, 50.86631, 57.9467, 58.74919,
    57.75268, 56.74033, 54.39473, 51.37042, 49.03791, 45.94575, 44.28364,
    42.99693, 40.73012, 39.00482, 31.63309, 22.97621, 18.86708, 17.85917,
    16.7491, 16.55237,
  60.24434, 53.43772, 47.15465, 47.89812, 57.2818, 62.62869, 63.52382,
    59.87384, 60.68097, 57.54737, 45.94577, 48.62531, 53.26463, 54.51313,
    52.47567, 51.90845, 49.72765, 43.73373, 40.76812, 38.99994, 38.07943,
    37.36811, 35.65342, 36.8292, 35.71412, 27.00803, 20.8499, 20.22386,
    18.10282, 16.70746,
  62.18307, 58.96511, 58.84978, 62.81398, 68.87691, 69.34106, 71.14305,
    66.74039, 65.87209, 55.79284, 44.98873, 52.39419, 56.29041, 58.12191,
    56.03682, 54.05138, 51.08424, 45.19355, 39.80926, 37.83515, 36.16586,
    34.50301, 33.45854, 32.87868, 33.85781, 33.22715, 27.4286, 21.69013,
    19.88092, 17.52424,
  64.86304, 66.97594, 62.65795, 65.80981, 70.30835, 69.6861, 67.07446,
    67.12436, 71.52589, 61.04625, 46.71701, 54.80272, 57.80841, 59.96283,
    58.30917, 56.77326, 51.94175, 46.81267, 41.58494, 37.05891, 36.37148,
    35.95185, 33.45743, 30.75964, 30.24602, 33.4854, 33.39569, 27.05689,
    23.97702, 20.40882,
  75.04333, 80.93224, 80.30471, 75.7672, 72.05531, 69.228, 73.27579,
    77.78711, 71.42151, 57.02507, 53.11349, 58.86175, 61.71872, 60.04044,
    55.86842, 54.38376, 50.72719, 46.74358, 42.99721, 38.56619, 37.41579,
    35.77962, 31.48697, 28.85853, 29.83125, 32.72176, 35.20446, 30.79343,
    23.3806, 20.08452,
  88.2086, 92.1162, 81.61074, 73.37449, 70.02054, 67.85828, 75.35757,
    75.99735, 62.69849, 53.66267, 58.59296, 61.63652, 61.21963, 57.8578,
    54.45062, 51.68538, 48.08715, 44.41994, 40.9059, 37.41964, 38.5762,
    41.31531, 40.47839, 37.5521, 37.65192, 39.3802, 42.1073, 37.70688,
    23.86431, 17.55968,
  93.60282, 87.97377, 77.061, 76.59208, 76.98852, 74.01332, 75.43225,
    68.77605, 55.71575, 57.25965, 60.36433, 60.71003, 59.12901, 56.50632,
    54.7822, 50.69912, 45.64347, 43.65194, 44.90256, 47.12629, 48.88412,
    47.6497, 43.12286, 41.02571, 41.07513, 42.97741, 44.06024, 45.2435,
    36.89291, 21.15127,
  79.15507, 73.30321, 78.47501, 86.50868, 86.74823, 85.43448, 77.22016,
    61.41271, 53.1924, 55.11286, 51.60624, 49.56789, 50.18848, 51.57062,
    53.56114, 54.01619, 53.58292, 54.09888, 51.62091, 47.47434, 45.70348,
    42.02762, 37.78983, 36.00089, 36.92752, 38.26185, 37.9369, 35.3581,
    32.35175, 24.36906,
  76.24689, 78.2878, 80.10905, 79.29976, 79.49329, 84.5643, 82.37152,
    63.45061, 51.70414, 55.53228, 56.83576, 60.12323, 63.03474, 63.9092,
    62.74924, 60.64094, 55.17086, 47.37184, 42.56411, 38.00678, 34.52689,
    32.67287, 31.11183, 30.23433, 30.3701, 31.02762, 30.13996, 25.94022,
    21.71853, 17.43098,
  23.9738, 24.31183, 24.8838, 25.6515, 26.32829, 27.34172, 28.56523,
    29.97963, 31.64996, 33.88175, 37.10978, 38.42738, 36.26715, 38.18385,
    39.57583, 39.41227, 40.07644, 41.44319, 42.99167, 45.30742, 46.57245,
    45.56484, 46.74909, 49.34745, 50.86817, 50.50894, 54.57294, 55.88927,
    38.69278, 32.52013,
  25.80204, 26.77639, 26.99349, 29.01435, 29.7879, 31.02161, 33.18575,
    35.43072, 37.93944, 40.79081, 44.25205, 48.0528, 50.63651, 50.34198,
    50.65528, 51.86266, 51.32008, 53.07932, 55.47717, 57.82584, 58.64871,
    58.73343, 59.21497, 62.14284, 64.62616, 58.07912, 50.15277, 53.72327,
    39.24112, 34.11682,
  28.75284, 30.57751, 32.56271, 34.70219, 36.64509, 38.59501, 40.47373,
    42.43978, 44.56305, 46.66676, 48.94135, 51.7049, 54.37074, 57.3288,
    59.33265, 57.97791, 59.40876, 62.45503, 65.7067, 71.07729, 78.78436,
    85.31044, 85.38596, 81.17769, 77.15541, 70.49277, 61.09297, 50.27103,
    37.86569, 34.62322,
  36.38554, 39.44082, 43.0083, 46.65945, 49.56437, 52.184, 53.13879,
    53.25795, 54.25785, 55.38644, 55.73161, 56.53489, 56.51954, 56.52748,
    60.63217, 62.92287, 60.51085, 59.06305, 64.54507, 71.13194, 80.43494,
    82.32195, 77.52013, 82.40282, 81.0493, 78.45502, 73.27004, 57.28429,
    41.79242, 33.21736,
  46.44761, 49.07039, 53.10851, 56.32892, 58.40625, 59.14628, 60.13769,
    60.99281, 63.1455, 64.85862, 64.97626, 67.37633, 68.71401, 68.57778,
    69.02837, 69.22139, 66.01489, 61.71593, 63.74072, 70.37705, 71.17119,
    63.06581, 65.50003, 72.93625, 79.35698, 79.75272, 74.61734, 79.66174,
    69.67601, 42.09531,
  61.31973, 67.23414, 71.83348, 75.73997, 74.56782, 73.34156, 75.85678,
    76.02567, 74.81107, 76.0508, 80.1447, 89.65312, 98.73177, 94.6377,
    93.69008, 93.52636, 90.58832, 82.23936, 71.94157, 70.36789, 62.90313,
    55.58526, 61.35532, 66.48899, 72.09109, 71.98752, 70.50572, 82.40901,
    72.59277, 37.69252,
  66.6832, 71.40291, 75.27263, 78.90276, 79.27464, 81.03093, 87.50414,
    91.98241, 88.99004, 82.79374, 77.61005, 69.00205, 59.11013, 60.83787,
    62.70972, 65.28424, 66.65017, 63.99044, 59.2241, 61.34391, 59.91331,
    59.53576, 63.53392, 68.87045, 69.54196, 64.39985, 67.78459, 74.58575,
    60.47441, 30.75848,
  59.73867, 64.04644, 69.41924, 74.22624, 76.56377, 84.0542, 87.36073,
    70.93694, 62.54715, 64.43356, 63.09076, 61.76194, 60.95618, 63.11997,
    64.5884, 67.00308, 69.55055, 68.03269, 63.15271, 63.88243, 65.12424,
    68.71113, 73.62956, 75.15736, 70.53812, 69.63148, 76.30043, 72.70573,
    51.26829, 32.58512,
  72.96796, 77.15514, 80.99591, 83.99048, 85.74889, 88.4458, 79.89632,
    80.88068, 86.09953, 89.32315, 91.327, 92.25114, 93.69469, 100.9556,
    102.9092, 88.90648, 86.2426, 86.67435, 83.30494, 76.83585, 73.86729,
    81.47824, 89.14469, 86.00667, 76.47285, 80.45875, 77.82993, 61.75864,
    35.64008, 32.07152,
  103.7734, 105.4148, 104.6209, 104.699, 104.3849, 98.45532, 80.50265,
    88.75269, 88.84082, 92.22025, 96.05149, 102.0372, 98.19942, 92.30721,
    87.30537, 91.32122, 91.5893, 88.5585, 83.93845, 83.61784, 85.78552,
    80.70114, 75.01892, 67.64963, 71.93755, 79.60329, 68.2901, 42.7709,
    31.34083, 29.40128,
  105.5916, 104.5471, 105.4036, 104.6574, 105.9299, 106.0001, 101.6299,
    103.0664, 102.5552, 94.96254, 78.49874, 59.7859, 56.52116, 56.59394,
    56.96497, 58.76764, 61.88306, 63.48435, 64.75763, 69.46405, 78.67404,
    73.30455, 59.66406, 57.62723, 62.26299, 58.33724, 42.07718, 32.37213,
    31.93441, 29.5829,
  111.2532, 107.1538, 109.4681, 109.4677, 108.5954, 105.4871, 100.4226,
    90.65276, 81.04914, 70.70841, 64.78947, 61.21333, 63.32418, 63.27071,
    59.55589, 57.35723, 55.61097, 56.10342, 57.49884, 62.87345, 71.73266,
    68.71516, 57.21313, 66.02481, 67.86684, 51.46041, 33.29345, 37.05991,
    33.38952, 31.02745,
  116.3146, 115.8632, 117.1721, 117.6002, 116.4344, 112.3179, 104.8233,
    101.1663, 102.6873, 99.81051, 94.01176, 87.16167, 92.17271, 92.63985,
    80.5536, 65.35235, 65.66679, 64.03892, 63.047, 67.34843, 68.45567,
    60.65723, 54.06131, 49.88663, 48.77192, 42.9217, 34.59963, 35.85589,
    35.15917, 32.2706,
  104.9212, 105.3297, 105.4956, 105.3122, 105.034, 105.3884, 106.0692,
    106.2496, 104.1949, 104.0901, 104.7362, 103.337, 104.2521, 104.5863,
    102.007, 82.94503, 77.88806, 81.61702, 83.45372, 75.37042, 63.34015,
    53.9959, 48.17146, 40.18142, 35.53011, 35.01874, 32.90375, 31.89369,
    32.32449, 31.5036,
  101.6393, 102.5005, 103.0539, 103.5917, 103.9559, 104.7139, 106.2581,
    105.6999, 103.6946, 103.4267, 95.77882, 89.5095, 90.78111, 92.63455,
    90.60205, 87.89755, 77.27129, 73.45916, 72.29637, 66.00185, 49.7886,
    48.68038, 41.28736, 38.25109, 37.01558, 35.25723, 33.49307, 31.93975,
    30.81411, 30.14519,
  104.1445, 105.3659, 105.5935, 105.3878, 105.0557, 105.5105, 106.1828,
    98.39051, 85.25798, 79.33427, 77.48087, 71.5268, 67.87371, 74.36121,
    71.26263, 68.59019, 68.78844, 61.46521, 59.58639, 53.61575, 41.9664,
    43.6817, 39.20539, 37.80392, 36.72551, 34.96103, 32.94009, 32.07526,
    31.11859, 30.24104,
  87.3148, 86.26503, 88.42556, 91.21873, 92.8066, 93.82602, 92.8189, 92.1131,
    88.9862, 82.2224, 74.74261, 82.938, 90.34124, 81.00116, 72.80952,
    65.5078, 58.94548, 56.34708, 57.61696, 53.38114, 41.67598, 43.62442,
    39.91006, 37.45953, 35.80843, 34.53601, 32.07014, 30.42514, 30.32358,
    30.01119,
  79.39713, 82.54948, 81.19887, 83.28928, 83.6965, 84.33258, 85.43771,
    85.35581, 85.35152, 85.40445, 94.60947, 103.0287, 99.56738, 96.5071,
    88.43187, 76.05574, 65.39603, 63.18759, 65.54221, 58.127, 43.47324,
    43.31248, 40.26772, 38.23722, 34.47582, 33.00716, 32.06062, 29.91631,
    29.84006, 29.63947,
  91.21339, 82.62043, 69.77288, 62.56698, 62.81844, 62.26424, 63.48443,
    65.46062, 66.4164, 69.47438, 75.67578, 73.80501, 65.41116, 70.10664,
    72.46042, 74.78858, 81.42934, 86.62568, 83.98788, 72.93694, 54.6299,
    46.72223, 41.47638, 38.24726, 34.43885, 32.43481, 31.57399, 30.27884,
    29.81751, 29.67087,
  83.77774, 73.90979, 61.67657, 54.88947, 56.50732, 58.07464, 59.75295,
    60.9437, 62.8084, 67.42913, 65.98017, 53.74492, 53.6932, 53.82066,
    53.72157, 54.57988, 59.87897, 67.0113, 70.88198, 70.64304, 64.67567,
    55.83503, 45.68787, 40.8878, 36.98602, 33.1503, 31.71171, 30.35904,
    29.74136, 29.66139,
  75.8128, 66.98175, 56.9481, 52.05212, 53.15322, 53.84051, 54.21682,
    53.72595, 54.78949, 56.38424, 50.26112, 41.95807, 46.34604, 46.40944,
    45.34815, 44.71433, 46.78557, 50.08852, 54.09777, 57.18938, 59.87674,
    60.92854, 54.33666, 46.65514, 40.39596, 34.84928, 31.89843, 30.52904,
    29.77003, 29.66139,
  75.00814, 66.05783, 59.19745, 54.76536, 54.37982, 51.35709, 50.84637,
    49.68536, 51.9529, 51.28459, 41.87358, 37.83075, 40.49176, 40.86573,
    40.23052, 40.64178, 41.30294, 43.03925, 46.20272, 48.86917, 51.37753,
    52.90299, 53.91458, 53.21188, 46.36819, 36.95117, 32.85319, 31.57501,
    30.03341, 29.61259,
  78.39011, 74.34984, 64.67972, 61.71629, 63.60009, 63.01112, 58.89427,
    53.25793, 52.57146, 49.02139, 41.70543, 43.0301, 44.44508, 45.16943,
    43.94581, 44.76226, 44.90934, 42.92731, 43.66625, 45.44963, 46.86139,
    47.62455, 47.76369, 50.01833, 50.90495, 43.12039, 35.99758, 34.10312,
    31.83332, 29.81533,
  85.86517, 82.60391, 78.95496, 77.08482, 77.27035, 73.56142, 74.97144,
    71.51862, 70.05556, 62.01045, 53.92062, 58.29008, 60.66533, 61.68112,
    59.52094, 57.9859, 55.8143, 52.36216, 49.4733, 49.16945, 48.58857,
    48.08844, 47.59094, 47.5389, 49.64975, 50.4011, 44.60838, 37.17696,
    34.53353, 31.09451,
  84.20953, 80.96288, 70.76814, 69.59624, 69.33858, 68.33379, 67.65208,
    70.27562, 74.08739, 64.75361, 54.67342, 59.22495, 61.6062, 62.97594,
    62.13883, 62.12002, 59.54096, 57.48541, 55.57197, 53.3725, 52.31725,
    50.65806, 47.70433, 45.96779, 47.26626, 50.52502, 50.78114, 42.92618,
    37.52599, 33.5449,
  92.09068, 88.07492, 81.17549, 73.83743, 70.41852, 68.23512, 72.12904,
    74.90739, 70.45729, 61.41282, 60.37307, 62.78692, 64.81043, 63.73837,
    61.56936, 61.86287, 61.66, 60.88606, 60.8073, 59.65614, 58.90936,
    57.23285, 53.28046, 50.41052, 51.02997, 52.30262, 53.13848, 45.59209,
    35.24661, 32.34764,
  93.56627, 87.50709, 77.35808, 71.34102, 67.47054, 64.57729, 68.37314,
    68.87025, 63.65448, 60.51811, 63.73692, 66.04962, 66.83434, 65.68848,
    63.63677, 62.01056, 61.38394, 61.70975, 62.54859, 62.65083, 63.61983,
    65.09305, 63.98149, 61.01011, 61.09644, 62.09675, 63.62165, 56.91957,
    39.65947, 30.58104,
  92.51145, 86.74121, 81.31044, 79.922, 78.14252, 73.04178, 70.62178,
    65.46375, 58.92554, 60.07696, 61.11746, 62.50878, 63.10886, 62.7498,
    62.06019, 59.71922, 57.50032, 57.5943, 59.58215, 60.81752, 58.96265,
    55.07764, 51.58763, 51.17392, 52.84832, 54.8615, 56.63864, 59.13255,
    51.7353, 35.08828,
  77.83102, 74.70604, 77.3509, 80.20422, 83.20036, 84.2691, 74.57848,
    60.69513, 54.23102, 54.28416, 51.7387, 50.72095, 50.90683, 51.4414,
    52.1032, 51.76044, 50.01032, 48.92494, 46.88289, 44.269, 43.42064,
    42.35191, 40.08692, 38.73568, 40.08167, 41.59392, 41.81753, 40.16085,
    40.26226, 35.96912,
  64.63849, 64.91776, 63.73008, 61.80607, 65.3403, 71.15182, 70.12227,
    56.38988, 49.01574, 52.27427, 53.8065, 54.82839, 54.42875, 52.87225,
    50.23835, 47.3522, 42.1692, 37.04042, 36.31183, 35.65054, 34.29427,
    34.85229, 34.99842, 35.05313, 35.74601, 37.02151, 37.27763, 34.7511,
    31.76681, 29.59312,
  41.286, 42.38273, 43.20126, 44.14241, 44.81895, 45.66768, 46.58546,
    47.4838, 48.45874, 49.53098, 50.93361, 51.15981, 49.1827, 49.3531,
    49.20737, 48.10632, 47.42242, 47.29308, 47.20432, 47.49719, 47.09073,
    45.19783, 45.24858, 47.04308, 48.02969, 46.79475, 48.59632, 50.31181,
    39.42563, 34.81827,
  47.51462, 48.65716, 48.72051, 49.96488, 50.09045, 50.47305, 51.45494,
    52.45771, 53.63317, 54.86068, 56.30928, 58.14022, 59.41024, 58.6185,
    58.078, 58.30545, 57.687, 58.49416, 59.52467, 60.37048, 59.95911,
    58.58026, 57.65117, 59.47862, 61.08527, 53.988, 46.14371, 48.93341,
    39.4973, 35.76186,
  50.57968, 51.57569, 52.09479, 52.57225, 52.72533, 52.88806, 53.05772,
    53.34711, 53.75859, 54.17767, 54.8047, 56.06385, 57.31785, 58.84859,
    59.92075, 58.90509, 59.80666, 62.07685, 64.73058, 68.59959, 74.43393,
    79.30323, 78.67778, 74.90097, 71.03256, 64.69206, 55.84462, 46.63354,
    38.11708, 36.09114,
  56.51192, 57.57231, 58.71922, 59.82064, 60.40187, 61.11783, 61.02669,
    60.38812, 60.32935, 60.34778, 59.83153, 59.60976, 58.54472, 57.42394,
    59.25007, 60.183, 57.9894, 56.83036, 60.73028, 65.61485, 72.36005,
    73.06232, 68.85606, 72.65908, 71.59412, 69.78381, 66.13515, 53.85128,
    41.47042, 35.43487,
  61.65749, 61.95871, 63.27686, 64.04242, 64.21346, 64.2926, 64.78645,
    65.0571, 66.42868, 67.56395, 68.00673, 69.99332, 70.58635, 69.27489,
    68.65788, 68.19875, 64.53783, 59.89616, 60.20278, 64.43157, 63.73294,
    56.16643, 57.23421, 62.93046, 68.55969, 69.75914, 67.10014, 72.54048,
    65.1666, 42.69203,
  65.87833, 69.04784, 71.62144, 73.70671, 72.54755, 72.1179, 74.56299,
    74.73891, 73.32554, 73.29601, 75.64792, 82.60374, 89.55036, 86.6543,
    86.60078, 87.37961, 84.0257, 76.3605, 67.17783, 65.10401, 58.16269,
    50.98687, 54.73514, 57.82465, 62.03098, 63.45197, 64.28329, 75.55815,
    68.92838, 38.825,
  71.34654, 75.41974, 78.47726, 81.10471, 81.59952, 83.91185, 89.58194,
    93.22832, 91.11462, 85.55717, 80.37321, 71.22874, 60.98948, 61.32918,
    62.07088, 63.8861, 64.65796, 61.28581, 57.39923, 58.02705, 55.9869,
    54.59059, 56.73951, 60.10983, 60.74776, 58.02805, 61.69743, 67.91997,
    56.13545, 33.25588,
  74.3085, 77.22763, 80.21031, 82.98161, 84.10881, 89.60397, 91.9825,
    78.28114, 71.85637, 72.15041, 69.40839, 66.3502, 63.83317, 63.53825,
    62.86148, 63.19601, 64.71097, 63.34827, 59.55495, 58.93248, 58.83714,
    60.68111, 63.90088, 65.53108, 63.02719, 62.98974, 68.1051, 65.16891,
    48.15887, 34.27696,
  79.94615, 79.75673, 79.61948, 79.90002, 80.32462, 80.65737, 71.41794,
    71.22464, 74.44809, 75.44256, 76.04537, 76.12251, 76.05093, 80.90398,
    82.47594, 74.19305, 73.05721, 73.83647, 71.84105, 66.42355, 63.01987,
    66.58398, 71.4784, 70.49437, 65.84138, 70.18723, 69.85616, 57.45935,
    36.4893, 34.34382,
  101.5578, 101.6587, 92.83354, 89.73343, 88.15144, 80.79846, 65.00998,
    69.31685, 67.68164, 68.25842, 69.58512, 73.72746, 73.23138, 70.90919,
    69.04688, 73.14098, 74.65995, 73.44965, 70.64757, 70.09871, 71.15047,
    67.7661, 63.41798, 58.70576, 62.68479, 70.26422, 62.58715, 42.0691,
    34.01834, 32.67739,
  108.4345, 107.564, 107.6948, 105.6707, 105.289, 94.78721, 85.31781,
    83.83826, 82.50162, 77.6633, 66.33505, 54.46678, 52.41757, 52.5271,
    52.79968, 54.17673, 56.12693, 57.23784, 57.98713, 60.70941, 67.354,
    64.99155, 56.10919, 55.24881, 58.92056, 55.49005, 42.20832, 34.58496,
    34.38994, 32.80467,
  114.7242, 111.7232, 113.213, 112.3734, 109.9326, 106.9604, 98.60443,
    88.62658, 81.2999, 74.24879, 68.51044, 64.06032, 64.37834, 62.74997,
    57.37711, 55.13266, 53.66645, 53.0266, 53.02667, 55.65473, 61.08097,
    59.74952, 52.97836, 59.47682, 62.05792, 49.53647, 35.41205, 38.07266,
    35.28478, 33.71442,
  110.7355, 111.6839, 112.6972, 113.2789, 113.0266, 110.6708, 105.1635,
    102.0648, 102.475, 94.74106, 89.14061, 82.80499, 85.88451, 85.67599,
    75.05814, 61.58154, 61.53592, 59.81655, 57.87992, 59.08244, 59.42988,
    54.52029, 49.87069, 46.23807, 46.10409, 42.23486, 36.48377, 37.13634,
    36.64411, 34.58897,
  93.08372, 93.683, 89.08042, 89.21723, 90.0332, 98.47013, 105.0393,
    104.7098, 94.37243, 97.74753, 102.1256, 98.55768, 97.98383, 97.43681,
    88.86559, 74.18137, 67.70165, 71.44025, 72.75772, 66.27723, 57.59123,
    50.20119, 45.47033, 39.67036, 36.54463, 36.47592, 35.17904, 34.38959,
    34.70045, 34.09985,
  75.24789, 71.85106, 73.27249, 73.44291, 74.38046, 76.24026, 80.57659,
    78.79599, 74.59584, 74.45712, 72.11316, 69.1746, 71.99192, 75.69357,
    74.63359, 73.67525, 67.51524, 64.1877, 63.08836, 58.5547, 47.87379,
    46.08399, 40.32738, 38.27816, 37.85753, 36.68343, 35.45367, 34.33976,
    33.53414, 33.11994,
  76.39887, 79.44578, 80.39874, 80.17276, 79.38548, 80.9947, 83.27298,
    78.80029, 72.21696, 68.71878, 67.53694, 63.98893, 61.96134, 64.91937,
    61.8736, 59.99871, 60.46783, 55.93444, 53.19548, 48.70019, 41.52599,
    41.7381, 38.77338, 37.954, 37.53175, 36.55514, 35.1136, 34.41511,
    33.69311, 33.13239,
  64.43863, 64.12704, 65.87224, 68.85306, 71.70148, 74.28818, 76.74485,
    79.36302, 78.11109, 74.28239, 70.36004, 75.71893, 80.00465, 73.75918,
    66.57902, 60.96016, 56.56082, 54.16291, 53.0681, 49.20791, 41.67188,
    42.15004, 39.35958, 37.79999, 37.01113, 36.34085, 34.60127, 33.33454,
    33.21524, 32.99262,
  55.96858, 56.15609, 55.58099, 58.23026, 61.23665, 64.48676, 67.03194,
    69.63441, 71.72084, 72.08635, 77.87578, 82.89114, 82.14104, 81.98846,
    77.63078, 71.01785, 65.24722, 63.08, 62.06739, 54.67979, 43.85118,
    42.29811, 40.01624, 38.58167, 36.36914, 35.42179, 34.57619, 33.02597,
    32.90574, 32.77244,
  61.69664, 55.80576, 48.632, 45.89083, 48.80119, 50.30618, 52.64069,
    55.01522, 55.88808, 58.38798, 62.22919, 61.16021, 57.394, 60.74767,
    62.61312, 64.91911, 70.99989, 75.53792, 73.60484, 65.2913, 52.37498,
    44.84482, 40.65954, 38.7095, 36.40108, 35.03582, 34.29306, 33.22667,
    32.88722, 32.8008,
  58.10502, 52.89007, 46.21958, 42.64801, 44.75855, 46.21383, 48.11775,
    49.96773, 52.48268, 56.81422, 56.85026, 50.67048, 50.92882, 50.17918,
    49.38718, 50.03641, 53.71803, 59.00345, 61.52201, 61.1813, 56.79875,
    50.25326, 43.51325, 40.39848, 37.98834, 35.53438, 34.41772, 33.34435,
    32.87508, 32.8117,
  60.02531, 55.35423, 48.11727, 44.66715, 45.38818, 45.95647, 47.11446,
    48.43736, 50.55059, 52.52298, 49.74522, 46.06014, 48.78657, 48.29809,
    46.7518, 45.97968, 46.99922, 48.8007, 50.49683, 50.91872, 51.66605,
    52.08887, 48.46748, 44.02532, 40.02196, 36.43956, 34.43647, 33.41078,
    32.89994, 32.80481,
  68.1974, 64.71201, 57.46448, 54.31161, 54.39683, 52.675, 52.71274, 52.6579,
    54.89388, 54.78276, 49.33278, 46.60637, 47.7612, 47.33006, 46.25446,
    45.87432, 45.38954, 45.63958, 46.56297, 46.83695, 47.13583, 47.32103,
    47.87915, 47.58936, 43.55869, 37.77213, 35.08109, 34.10596, 33.10341,
    32.80497,
  73.63927, 73.82199, 66.41923, 64.68943, 66.76147, 67.01039, 65.11051,
    61.63989, 61.5256, 59.54913, 54.70758, 54.8191, 54.60963, 53.68148,
    51.60517, 51.05081, 49.84824, 47.24924, 46.35272, 45.86602, 45.25014,
    44.75189, 44.47574, 45.78699, 46.6359, 41.95419, 37.26715, 35.91504,
    34.37167, 32.95987,
  75.89252, 75.74213, 71.78436, 70.98876, 71.89964, 71.80122, 72.39465,
    71.48586, 72.99765, 68.11484, 63.26283, 65.40088, 65.91729, 65.32328,
    62.91542, 60.83891, 58.12642, 54.43729, 51.16261, 49.11303, 47.20938,
    45.8092, 45.04568, 44.78495, 46.22694, 46.7259, 42.88021, 38.05772,
    36.21807, 33.80556,
  76.75241, 72.83829, 66.81883, 65.18707, 65.94984, 65.92675, 67.35389,
    71.18053, 75.27456, 70.07977, 63.57943, 65.41962, 66.05817, 66.38431,
    65.15118, 63.84595, 60.67575, 57.80143, 55.19648, 52.48564, 50.54532,
    48.30426, 45.57327, 43.89953, 44.85286, 47.10564, 47.23235, 41.81472,
    38.1664, 35.37965,
  79.59167, 76.20045, 70.27442, 65.71329, 63.66808, 63.1505, 67.08316,
    71.50151, 70.63833, 65.57296, 65.04385, 65.74948, 66.39862, 65.37273,
    63.25708, 62.39786, 61.06914, 59.46927, 58.5128, 56.61938, 55.64664,
    53.92319, 49.89448, 46.71861, 46.76467, 47.81162, 48.67823, 43.64173,
    36.61214, 34.46949,
  77.09711, 72.86039, 65.99901, 62.38086, 59.83233, 57.1889, 60.2121,
    61.6362, 59.70725, 58.14269, 60.14591, 61.59759, 62.1664, 61.96307,
    60.7291, 59.43366, 58.23445, 57.85527, 57.7587, 57.02666, 57.26689,
    57.99707, 56.30404, 53.30445, 52.56132, 53.52265, 54.95137, 50.60435,
    39.47512, 33.42566,
  70.0229, 68.17259, 64.63544, 63.05447, 62.43627, 59.24369, 56.74657,
    53.63305, 50.20959, 50.904, 51.88526, 53.55341, 55.09001, 55.95024,
    56.15598, 55.12621, 53.36208, 52.8601, 53.8141, 54.26291, 53.15295,
    50.68069, 47.87986, 47.19439, 48.04314, 49.16492, 50.2753, 51.78688,
    47.00323, 36.34592,
  55.38548, 55.10493, 56.30272, 57.47349, 59.68799, 61.5144, 56.35094,
    47.93827, 45.37207, 46.73895, 46.47106, 46.65722, 47.41428, 47.87344,
    48.19021, 48.21969, 46.93724, 45.87248, 44.53469, 42.85041, 42.35131,
    41.70547, 40.24514, 39.44007, 40.25446, 40.85659, 40.63754, 39.59943,
    39.66187, 36.81757,
  45.6919, 46.34902, 45.96641, 44.98985, 47.08385, 51.72084, 52.29681,
    44.74471, 40.98529, 43.50315, 45.10963, 46.50299, 46.89668, 46.02578,
    44.60656, 43.52054, 40.54837, 37.38327, 37.09361, 36.7064, 35.83924,
    36.29001, 36.57185, 36.66005, 37.02143, 37.67889, 37.62742, 36.16191,
    34.39497, 32.81705,
  44.75991, 44.86816, 44.98945, 45.18304, 45.12805, 45.18245, 45.27599,
    45.42215, 45.72997, 46.31734, 47.31496, 47.27087, 45.51472, 46.08273,
    46.46222, 46.22703, 46.63728, 47.50008, 48.36485, 49.52071, 49.7901,
    48.45875, 48.83638, 50.54506, 51.69408, 51.19524, 52.73516, 53.90918,
    44.63357, 41.244,
  48.85078, 49.20401, 48.82403, 49.49299, 49.2701, 49.27983, 49.75891,
    50.17416, 50.77493, 51.59309, 52.56868, 53.77832, 54.59511, 53.96083,
    53.71989, 54.338, 54.18534, 55.32253, 56.77085, 57.93789, 57.98475,
    57.49661, 57.62821, 59.98986, 62.19937, 57.12372, 49.85862, 53.00215,
    44.88412, 41.99373,
  49.67437, 49.95596, 50.13329, 50.38237, 50.62085, 51.00512, 51.54523,
    52.27213, 53.17332, 54.14055, 55.23171, 56.76042, 58.32637, 60.14749,
    61.45199, 60.65067, 61.75598, 63.88706, 66.11256, 69.30931, 74.556,
    79.56956, 78.80138, 73.7539, 69.95291, 65.4375, 58.52096, 51.39436,
    44.28964, 42.52952,
  53.33089, 53.68702, 54.25275, 54.93415, 55.3474, 55.90112, 56.07854,
    56.06348, 56.59599, 57.22902, 57.53045, 58.29354, 58.7051, 58.87937,
    61.46595, 63.19493, 62.24121, 62.08656, 65.68385, 70.03767, 76.20125,
    76.37658, 70.56174, 72.15756, 69.60452, 68.26786, 66.6693, 55.71298,
    45.67648, 41.6522,
  58.47523, 58.40322, 59.2947, 59.80237, 59.94395, 59.89725, 60.3822,
    60.71603, 61.86871, 62.78159, 63.15902, 65.1106, 66.50092, 66.36656,
    67.04833, 68.30063, 67.16124, 64.62392, 66.08917, 70.69998, 70.59568,
    62.42884, 62.44881, 66.60431, 69.90401, 70.34038, 68.32859, 72.81725,
    67.30207, 49.01929,
  62.70997, 64.68592, 66.54948, 68.24445, 67.5797, 67.63967, 70.14768,
    70.94267, 70.65118, 71.48019, 74.43198, 82.01717, 89.53471, 87.24107,
    87.90113, 89.40447, 87.65821, 81.35344, 73.23369, 70.64276, 64.01026,
    56.96405, 60.9922, 63.91404, 67.57581, 68.70842, 69.72311, 79.38564,
    73.21257, 45.5309,
  63.98613, 66.31857, 68.48161, 70.60722, 71.25148, 73.59978, 79.64362,
    84.23854, 83.51808, 79.55171, 75.81732, 69.08285, 60.81089, 62.17572,
    63.89283, 66.10146, 67.27504, 65.21916, 61.67415, 61.53239, 58.83592,
    57.4559, 59.95931, 63.51051, 64.74284, 63.33416, 67.74834, 73.92276,
    62.29565, 39.98769,
  64.47113, 66.94375, 69.61813, 72.08097, 73.09978, 77.84709, 80.1166,
    68.02886, 62.31429, 63.11088, 61.41122, 59.52114, 58.39088, 59.25174,
    60.2883, 62.43504, 65.29002, 65.26328, 62.07339, 61.30447, 60.86242,
    61.83318, 64.42513, 66.2832, 65.3699, 66.64133, 72.6758, 70.46202,
    54.53741, 40.59245,
  70.33614, 71.5865, 72.67176, 74.00024, 75.61971, 76.22444, 67.58826,
    67.03049, 69.72937, 70.81747, 71.54964, 71.8675, 72.80542, 77.40273,
    79.42568, 73.54184, 74.42208, 76.39761, 74.69826, 69.82509, 66.92258,
    69.84606, 73.45562, 72.29614, 69.02641, 73.79931, 74.08015, 62.56206,
    42.74754, 41.16023,
  85.99677, 86.89956, 80.55171, 79.76657, 80.8279, 75.21936, 60.83983,
    66.06544, 65.85976, 67.59882, 69.96844, 74.46457, 74.52847, 73.26002,
    71.88091, 75.46742, 77.1004, 76.74398, 74.52576, 73.99933, 74.56982,
    71.50667, 68.40044, 64.64184, 69.02722, 76.18518, 68.24564, 48.54123,
    40.58048, 39.71927,
  99.17963, 98.18713, 98.04525, 90.80876, 90.91797, 81.2511, 72.5659,
    73.56848, 73.8821, 70.87511, 63.25157, 55.05673, 54.70587, 55.88621,
    56.64926, 58.38271, 60.65498, 61.93341, 62.69901, 65.40515, 70.9651,
    69.10174, 61.83365, 60.92953, 65.24567, 62.83334, 49.5029, 40.77114,
    41.14948, 39.7304,
  106.2877, 103.012, 104.2094, 103.0029, 100.3149, 90.23051, 83.86307,
    75.28485, 69.39436, 65.2393, 61.36153, 59.27848, 60.73425, 60.20332,
    57.7767, 57.14193, 57.05533, 57.63256, 58.30564, 61.11264, 66.3724,
    66.15175, 61.43329, 67.64581, 69.6434, 56.33572, 41.73717, 44.29144,
    41.73308, 40.46027,
  105.7558, 106.1979, 106.8497, 106.3835, 104.737, 101.5267, 95.34957,
    88.60178, 92.26509, 84.39174, 79.42889, 74.76019, 78.18822, 78.8336,
    71.65654, 61.47155, 62.0946, 61.9156, 61.19, 62.89853, 64.49376,
    61.97483, 58.71829, 55.75658, 54.78641, 49.84837, 43.18548, 44.0165,
    43.17935, 41.30413,
  95.35703, 96.35945, 93.80763, 93.12468, 92.26934, 94.20173, 94.54385,
    94.34261, 91.32632, 92.4612, 92.25928, 91.07188, 91.25031, 91.37886,
    88.05514, 73.77643, 70.45442, 73.60754, 75.73042, 69.65474, 61.96189,
    56.36992, 52.17297, 46.39223, 43.57289, 43.34978, 42.14948, 41.45853,
    41.54646, 40.93081,
  69.64392, 66.01722, 67.96286, 68.39902, 69.8847, 72.23303, 76.3765,
    76.17403, 73.21222, 73.85328, 72.39005, 70.21985, 73.90994, 78.89514,
    79.57379, 77.63546, 70.48567, 67.75784, 66.12188, 62.26843, 53.2269,
    51.40504, 46.29931, 44.1909, 44.00415, 43.19284, 42.07032, 41.10174,
    40.40075, 40.04718,
  68.62538, 70.36375, 70.64757, 70.12697, 69.14299, 70.11325, 71.96222,
    69.51435, 65.20935, 63.11673, 63.03954, 61.41818, 61.35976, 65.05623,
    63.28397, 62.20545, 63.02771, 59.03392, 56.81779, 52.89367, 47.02922,
    47.22727, 44.65007, 43.88001, 43.83044, 43.19452, 41.90816, 41.18367,
    40.51114, 40.03875,
  62.1026, 61.43711, 62.20864, 63.87769, 65.46527, 66.65471, 67.84705,
    69.51471, 68.57133, 66.13447, 62.86124, 67.2804, 72.10771, 68.19105,
    62.74153, 59.42205, 57.17913, 56.01208, 55.70665, 53.10406, 47.20042,
    47.49101, 44.96116, 43.76068, 43.50745, 43.13506, 41.62507, 40.42045,
    40.19139, 39.97947,
  56.99147, 57.7605, 57.17947, 59.13157, 61.17764, 63.28684, 64.91518,
    66.58972, 67.98773, 67.85594, 71.759, 75.30891, 75.14579, 74.86438,
    70.6669, 65.96146, 61.39783, 60.43665, 60.52128, 55.69127, 48.19345,
    47.38482, 45.48353, 44.55173, 43.08384, 42.29192, 41.45992, 40.08031,
    39.92758, 39.78275,
  63.31452, 58.89644, 52.6591, 50.04721, 52.55127, 53.70457, 55.56709,
    57.51805, 58.43486, 60.7906, 64.58223, 64.33236, 61.07479, 63.42117,
    64.42348, 66.45928, 71.26328, 74.81331, 72.61964, 65.42582, 55.0253,
    49.24357, 46.01337, 44.77505, 43.06748, 41.90124, 41.20943, 40.19919,
    39.88938, 39.79602,
  60.10214, 55.69034, 49.44144, 46.01262, 47.67821, 48.65696, 50.03552,
    51.5834, 53.80236, 57.45129, 58.35357, 54.56083, 55.31012, 55.07374,
    54.78669, 55.62762, 58.83193, 63.05809, 64.16998, 62.70316, 58.1945,
    52.74361, 47.95706, 46.09634, 44.41863, 42.27171, 41.3043, 40.32101,
    39.88133, 39.81607,
  59.09385, 54.70364, 48.05591, 44.64974, 45.26299, 45.72232, 46.66209,
    47.91434, 49.94561, 52.03759, 50.67984, 48.46728, 51.36475, 51.76729,
    51.06575, 51.03299, 52.22456, 53.7429, 54.96476, 54.79675, 54.69922,
    54.37753, 51.43948, 48.60505, 45.75335, 42.91587, 41.27388, 40.31609,
    39.8631, 39.79789,
  62.64663, 59.00635, 52.25846, 48.95462, 49.05728, 47.93563, 48.32677,
    48.71432, 50.98271, 51.52611, 47.92908, 46.69095, 48.59935, 49.11769,
    48.94007, 49.40865, 49.71612, 50.36002, 51.30822, 51.76408, 51.91427,
    51.75917, 51.83181, 51.10655, 47.90383, 43.51928, 41.61295, 40.74604,
    39.95287, 39.7693,
  67.86031, 66.84774, 59.20873, 56.60827, 58.0145, 58.06448, 56.84734,
    54.63335, 54.75328, 53.5028, 50.09497, 50.93028, 51.83324, 52.11,
    51.32808, 51.8302, 51.8732, 50.48582, 50.19276, 50.11506, 49.7612,
    49.3275, 48.947, 49.62398, 49.81973, 46.06219, 42.9644, 41.98322,
    40.83178, 39.88,
  71.38213, 70.93845, 65.94865, 64.23225, 64.7513, 64.18433, 64.75962,
    64.33831, 65.71509, 62.58271, 58.85724, 61.12866, 62.5499, 62.76833,
    61.23149, 60.182, 59.13487, 56.92807, 54.27679, 52.66553, 51.33015,
    50.49745, 49.67272, 49.22805, 50.11891, 50.21898, 47.20938, 43.35068,
    42.06726, 40.4859,
  71.64896, 68.15157, 62.70591, 60.7572, 61.45976, 61.33265, 62.34342,
    65.1817, 68.50809, 65.0415, 60.42984, 62.35168, 63.87439, 64.76221,
    63.86352, 63.37944, 62.44909, 61.01165, 58.32308, 55.84279, 54.36487,
    52.62645, 50.30087, 48.99673, 49.79748, 51.47481, 51.19893, 46.63549,
    43.82318, 41.74157,
  73.10081, 70.31194, 65.62225, 62.01808, 61.3102, 61.32959, 64.71705,
    68.37453, 67.72784, 63.4763, 63.22033, 64.30114, 65.62216, 65.2982,
    63.57485, 63.28346, 63.4874, 62.78386, 60.78313, 58.56281, 57.80958,
    56.28628, 52.81483, 50.57837, 50.86697, 51.53883, 51.91652, 48.11124,
    42.81628, 41.18835,
  72.04785, 68.86978, 64.15456, 61.26237, 60.13487, 59.03234, 62.21498,
    63.88491, 62.79319, 61.60754, 63.41318, 64.80853, 65.75135, 65.73963,
    64.70072, 64.04762, 64.19858, 64.08607, 62.59292, 61.20718, 61.66926,
    62.09653, 60.15853, 57.51447, 56.60165, 56.52665, 56.67043, 52.79068,
    44.29613, 40.24448,
  66.99162, 65.01415, 62.36465, 61.94649, 61.98876, 60.38247, 59.45634,
    57.87233, 55.71774, 56.77439, 58.23093, 60.04788, 61.75594, 62.86837,
    63.08083, 62.6747, 62.04591, 61.65524, 61.33748, 61.07031, 60.08017,
    58.0428, 55.51694, 54.5825, 54.88841, 55.09578, 54.80877, 55.01167,
    50.73697, 42.41227,
  56.02738, 56.15931, 57.06059, 58.01482, 60.03775, 61.78587, 58.43816,
    52.22256, 50.41756, 51.36447, 51.19486, 51.79915, 53.11597, 54.48597,
    55.50284, 55.82447, 55.13602, 54.15448, 52.39861, 50.54962, 49.84019,
    49.14367, 47.90572, 47.17873, 47.76516, 48.10035, 47.44793, 46.11166,
    45.84784, 43.30608,
  50.43659, 51.16148, 51.18443, 50.67597, 52.60036, 56.74256, 57.42879,
    51.29277, 48.43134, 50.47495, 51.82313, 53.30085, 53.78973, 53.19196,
    51.75092, 50.45362, 48.02184, 45.75611, 45.30224, 44.62355, 43.74313,
    44.06176, 44.41988, 44.41359, 44.62213, 44.80054, 44.27863, 42.84415,
    41.39069, 39.91589,
  42.75664, 42.88399, 43.0566, 43.22438, 43.34714, 43.57535, 43.839,
    44.13876, 44.51104, 45.08804, 45.96337, 45.75639, 44.08465, 44.4707,
    44.6291, 44.30937, 44.4633, 44.85197, 45.38631, 46.32073, 46.92752,
    46.52872, 47.14502, 48.9208, 50.55124, 50.69329, 52.18028, 53.36484,
    46.20913, 43.65902,
  45.15134, 45.44367, 45.19948, 45.7286, 45.61891, 45.65262, 45.91751,
    46.17999, 46.53774, 46.96678, 47.51423, 48.08274, 48.35848, 47.59381,
    47.28681, 47.83812, 47.67061, 48.53154, 49.65684, 50.86847, 51.57325,
    52.22916, 53.96161, 58.03719, 61.42025, 56.77368, 50.04257, 52.98642,
    46.5703, 44.26507,
  47.30654, 47.68498, 47.96074, 48.23946, 48.4193, 48.6817, 48.97109,
    49.35214, 49.83762, 50.34621, 50.95041, 51.87696, 52.95329, 54.33287,
    55.32212, 54.95808, 56.21875, 58.03174, 60.01482, 63.04805, 68.12165,
    73.89597, 75.03225, 71.73063, 68.80246, 63.53185, 58.00765, 51.79075,
    46.39442, 44.76628,
  51.53016, 52.42349, 53.39675, 54.39713, 54.9234, 55.48962, 55.62469,
    55.5935, 55.95585, 56.53598, 56.98989, 57.94186, 58.57358, 58.75637,
    60.92172, 62.36195, 61.79044, 61.94895, 64.93005, 68.79556, 74.64299,
    74.89119, 69.02981, 69.51904, 66.53932, 65.39758, 63.83651, 54.59561,
    46.48977, 43.81141,
  54.13829, 54.10158, 55.06537, 55.68088, 55.88107, 55.87623, 56.24461,
    56.48336, 57.26286, 57.6483, 57.78095, 59.14327, 60.35171, 60.95886,
    62.05178, 63.70701, 63.6707, 62.65604, 65.20766, 69.94669, 70.10495,
    62.29388, 61.17699, 64.97137, 67.60172, 67.82503, 66.85635, 71.49107,
    67.53407, 51.06179,
  57.73938, 59.53831, 61.40411, 63.21223, 63.27386, 64.03622, 66.83289,
    68.56031, 70.08184, 72.6053, 76.81069, 85.3856, 86.17755, 85.74334,
    85.9749, 86.41727, 85.75385, 81.88738, 75.11506, 72.50812, 66.27332,
    59.02365, 63.03485, 65.86444, 69.33772, 70.69538, 71.99276, 80.61984,
    74.40058, 48.38107,
  66.06867, 69.42732, 72.2289, 75.06496, 76.97385, 80.84026, 86.34995,
    86.53826, 86.20934, 85.76601, 85.47341, 81.22269, 72.98028, 73.24059,
    73.655, 74.26538, 74.25999, 70.08557, 65.46312, 64.42635, 60.95122,
    59.34542, 61.99246, 65.14037, 66.32797, 65.24072, 69.1823, 74.53722,
    63.25475, 42.57582,
  67.72054, 70.46478, 72.83074, 75.28228, 76.66869, 81.44527, 83.51718,
    71.45576, 64.81277, 64.27811, 61.54327, 58.72131, 57.06047, 57.83909,
    59.03466, 61.24201, 63.1062, 62.51149, 60.11092, 59.74255, 59.36491,
    60.40141, 63.18563, 65.48564, 65.25742, 66.91225, 72.94623, 71.34053,
    56.36569, 42.67783,
  68.20522, 69.63044, 70.75025, 71.80219, 73.73685, 74.05286, 65.23213,
    63.17792, 65.14727, 65.70798, 65.99954, 66.04568, 67.2273, 71.59673,
    73.67669, 69.2795, 70.68782, 72.63987, 71.45952, 67.56441, 65.56406,
    68.56853, 72.12233, 71.39722, 68.98335, 74.2917, 76.09152, 64.85846,
    45.2781, 43.52768,
  75.69763, 79.2296, 76.84142, 78.66316, 80.9727, 77.03867, 64.18956,
    69.80429, 70.98483, 74.01956, 76.97691, 80.11749, 79.2645, 77.58651,
    75.79347, 77.62527, 78.45578, 77.97263, 75.97003, 74.76419, 74.73219,
    72.34695, 69.58135, 66.36079, 70.11175, 77.24941, 70.83811, 51.19336,
    42.87743, 42.50925,
  81.4193, 81.77931, 83.23325, 83.15311, 86.66022, 81.10295, 73.96331,
    77.18433, 79.84932, 78.53889, 70.97927, 62.37185, 61.20011, 61.87025,
    62.17147, 62.83407, 64.03926, 64.59982, 64.86493, 66.76997, 70.83694,
    68.63162, 62.30113, 61.84357, 66.71551, 65.3652, 52.38608, 42.92422,
    43.56179, 42.4279,
  91.28462, 89.30506, 91.63279, 91.79114, 90.64091, 80.33757, 79.71621,
    72.16029, 66.65735, 65.46503, 61.46729, 59.31359, 60.96704, 60.92773,
    58.97251, 59.0604, 58.54729, 59.18251, 59.59979, 61.60535, 65.97156,
    65.85829, 62.05112, 67.46547, 69.28242, 57.70951, 43.703, 45.92839,
    43.95711, 43.0204,
  98.27831, 99.10571, 99.9642, 99.19434, 96.90109, 93.10467, 87.2039,
    80.23474, 85.34648, 77.47618, 73.42156, 70.34564, 74.0546, 75.32448,
    69.55547, 59.99249, 61.44521, 61.55356, 61.37736, 63.47237, 65.98613,
    65.20503, 62.55434, 59.15014, 57.05011, 51.91255, 45.25411, 46.20702,
    45.21598, 43.7929,
  93.6023, 93.47729, 92.64848, 90.45454, 88.97196, 88.68967, 88.75199,
    88.31257, 86.64571, 86.67647, 86.75369, 85.78893, 86.29376, 86.65192,
    85.31374, 74.02731, 70.07955, 74.60001, 76.17586, 70.40711, 64.47294,
    59.47018, 54.60098, 48.78772, 46.11006, 45.7313, 44.76509, 44.12826,
    44.08363, 43.52893,
  87.98087, 84.62691, 85.22246, 84.38353, 85.06323, 87.06639, 88.76897,
    88.40277, 86.03739, 85.30673, 82.30352, 79.12479, 79.75014, 82.20148,
    81.61047, 79.46599, 74.24253, 71.03907, 69.09372, 64.5218, 55.4133,
    53.0172, 48.05774, 45.61264, 45.63119, 45.31847, 44.50616, 43.61749,
    43.0539, 42.74507,
  74.43892, 75.79655, 76.21304, 75.4706, 74.28787, 75.29728, 76.90385, 74.56,
    70.45296, 68.0958, 67.8123, 65.91895, 65.5078, 68.63823, 66.58781,
    65.69357, 65.51152, 61.5403, 58.89628, 54.65845, 49.10592, 48.76679,
    46.09841, 45.41566, 45.47428, 45.27639, 44.45396, 43.73765, 43.14117,
    42.71897,
  64.23256, 63.23799, 63.56949, 64.33649, 65.13244, 65.65178, 66.57027,
    67.8048, 66.80542, 64.73074, 61.92803, 65.63885, 69.90292, 67.12521,
    62.63857, 60.17519, 58.30851, 57.0431, 56.60043, 54.12011, 48.73038,
    49.01721, 46.61089, 45.53304, 45.45536, 45.32725, 44.22821, 43.19158,
    42.92526, 42.7003,
  59.9712, 60.73431, 60.22437, 61.35588, 62.24324, 63.5358, 64.55775,
    65.56065, 66.37063, 65.73087, 68.54912, 71.33027, 70.72046, 69.65633,
    65.43884, 61.78409, 58.22689, 57.76939, 58.50616, 55.15915, 49.10083,
    48.75063, 46.95605, 46.22233, 45.21252, 44.67537, 44.02697, 42.85139,
    42.68523, 42.52049,
  69.62027, 65.3859, 59.37709, 56.51461, 58.02158, 58.24206, 59.22998,
    60.40203, 60.57611, 62.05137, 64.95767, 64.45911, 60.90773, 61.97689,
    61.79495, 63.2664, 67.49609, 70.8791, 69.3971, 63.27213, 54.7371,
    50.2088, 47.53369, 46.64088, 45.41373, 44.50264, 43.86637, 42.96185,
    42.66897, 42.55042,
  68.03706, 63.71185, 57.97068, 54.54469, 55.85172, 56.38757, 57.37466,
    58.45511, 60.07922, 62.7979, 63.35174, 60.02957, 59.99785, 59.2993,
    58.70636, 59.17554, 61.49828, 64.69801, 64.62941, 62.29717, 58.14351,
    53.21032, 49.10342, 47.8065, 46.53867, 44.8394, 43.92619, 43.0344,
    42.64474, 42.54113,
  65.00006, 61.37394, 55.73238, 52.6874, 53.62879, 54.08766, 54.88942,
    55.88401, 57.23351, 58.54678, 57.15642, 54.8944, 56.76522, 56.58384,
    55.54732, 55.07277, 55.47477, 56.13612, 56.5114, 55.58411, 55.12963,
    54.64274, 52.01117, 49.76228, 47.80561, 45.42828, 43.94611, 43.02975,
    42.62413, 42.54035,
  63.58052, 60.59719, 55.0463, 52.39787, 52.97583, 52.42288, 53.25843,
    53.90461, 55.67341, 55.88586, 52.73956, 51.3066, 52.62636, 52.77565,
    52.49761, 52.55587, 52.44129, 52.74997, 53.30452, 53.5391, 53.5693,
    53.2056, 52.91714, 51.79492, 49.1349, 45.77662, 44.17578, 43.3551,
    42.67849, 42.51783,
  63.15152, 61.62178, 55.52387, 53.51522, 55.06153, 55.3141, 54.72655,
    53.46741, 53.89232, 53.06248, 50.28252, 50.78544, 51.56716, 52.12226,
    51.84498, 52.46721, 52.62924, 51.76088, 51.6214, 51.52238, 51.3853,
    51.02861, 50.48457, 50.52517, 50.42046, 47.5494, 45.23931, 44.45803,
    43.44492, 42.61067,
  67.95995, 67.45523, 62.9941, 61.60642, 61.96966, 61.25399, 61.74833,
    61.52254, 63.0282, 61.15053, 58.43602, 59.99676, 61.08048, 61.39437,
    60.11144, 59.25422, 58.55095, 56.9077, 54.71424, 53.35861, 52.44304,
    51.89571, 50.99141, 50.36171, 50.78533, 50.67939, 48.32493, 45.38503,
    44.31405, 43.11586,
  71.13167, 68.45882, 62.71442, 60.62504, 60.91259, 60.59094, 61.59193,
    64.21198, 67.6395, 65.3729, 61.84859, 63.7992, 65.23737, 65.67709,
    64.22483, 63.70358, 63.09846, 61.7939, 59.37069, 56.97462, 55.50578,
    54.06874, 51.91794, 50.61474, 51.2065, 52.38323, 51.78768, 47.89063,
    45.69456, 44.17906,
  73.05115, 71.48295, 66.47379, 62.62732, 61.97369, 61.83083, 64.62258,
    68.23276, 68.51723, 64.6618, 64.29047, 65.59114, 66.78552, 66.02078,
    64.05988, 63.76067, 63.41275, 62.13522, 59.97849, 57.73852, 56.78461,
    55.44402, 52.65415, 51.03461, 51.5478, 52.11216, 52.29601, 49.09274,
    45.01266, 43.77834,
  74.30372, 71.88039, 67.29224, 64.13866, 63.20157, 62.15969, 64.8601,
    66.58762, 65.47794, 63.74118, 64.68132, 65.82161, 66.6507, 66.04504,
    64.68443, 63.92967, 63.40848, 62.4571, 60.93501, 59.85855, 59.99641,
    60.16469, 58.311, 56.15137, 55.62, 55.59, 55.58699, 52.32811, 45.87936,
    42.89068,
  74.23812, 72.5163, 69.30836, 68.71353, 69.20695, 68.09985, 67.61859,
    66.51243, 64.34523, 64.49107, 65.48529, 66.97428, 68.21216, 68.54525,
    68.00706, 67.05122, 65.71612, 64.83542, 64.55079, 64.30614, 62.92274,
    60.32835, 57.44189, 56.11143, 55.92296, 55.8915, 55.30741, 55.00861,
    51.34708, 44.5136,
  64.42415, 64.39699, 65.05104, 65.86461, 67.86149, 69.51872, 66.38701,
    60.88516, 59.21079, 59.68673, 59.3321, 59.70761, 60.74748, 61.90445,
    62.90358, 62.80804, 61.4015, 59.97193, 58.03104, 55.96402, 54.7106,
    53.35238, 51.65109, 50.58921, 50.71101, 50.70343, 49.90954, 48.59983,
    48.06146, 45.55315,
  59.95444, 60.28253, 60.41213, 60.1889, 62.33273, 66.14362, 66.21956,
    60.27717, 57.47477, 58.84194, 59.4872, 59.94573, 59.52978, 58.53791,
    57.36307, 56.0514, 53.36482, 50.95059, 50.10852, 49.0435, 47.95064,
    47.9502, 47.97648, 47.87573, 47.81074, 47.66523, 46.76061, 45.41234,
    44.21327, 42.75978,
  41.45452, 41.42722, 41.50342, 41.57566, 41.61375, 41.64645, 41.77816,
    41.99321, 42.28773, 42.71646, 43.3987, 43.20062, 41.97737, 42.34428,
    42.42263, 42.03935, 42.08076, 42.18813, 42.37202, 42.90239, 43.19076,
    42.76049, 43.11685, 44.4303, 45.86758, 46.24087, 47.61003, 48.99994,
    44.32172, 42.29269,
  42.3555, 42.423, 42.26997, 42.5653, 42.46787, 42.45583, 42.66367, 42.92921,
    43.24868, 43.61875, 43.98088, 44.23086, 44.28447, 43.57957, 43.09509,
    43.24097, 42.83143, 43.16454, 43.71437, 44.33084, 44.72623, 45.51047,
    47.80039, 52.41387, 56.39243, 52.56823, 46.81699, 49.5574, 44.85157,
    42.83575,
  42.51434, 42.42014, 42.43128, 42.44474, 42.43694, 42.58055, 42.75193,
    42.99355, 43.28656, 43.55707, 43.89053, 44.41402, 44.99501, 45.71848,
    46.15549, 45.76846, 46.68449, 48.24917, 50.15961, 53.33691, 59.03327,
    66.04085, 68.64624, 66.51021, 63.75343, 58.56886, 54.19824, 48.87938,
    44.66691, 43.26615,
  43.47576, 43.79194, 44.49121, 45.24643, 45.85244, 46.57255, 46.93694,
    47.0746, 47.41316, 47.94652, 48.36157, 49.2943, 50.00694, 50.37288,
    52.47869, 54.29886, 54.8897, 56.28895, 60.20396, 65.39054, 72.33749,
    72.76296, 66.43556, 65.3822, 61.38918, 60.48267, 59.65041, 51.40356,
    44.02337, 42.24601,
  46.75962, 47.06115, 48.07454, 48.81305, 49.06517, 49.17268, 49.33678,
    49.21058, 49.35497, 49.19854, 49.07841, 50.25559, 51.90954, 53.6797,
    55.83703, 58.36613, 59.61682, 60.33955, 63.78831, 68.64024, 68.38602,
    59.86121, 56.61534, 59.60653, 61.15488, 61.36296, 61.66953, 66.93781,
    64.25504, 49.38625,
  48.26361, 48.83154, 49.67971, 50.30817, 49.57441, 49.41626, 50.96365,
    52.49624, 54.66488, 58.12353, 63.59729, 73.6837, 82.82841, 82.23529,
    84.17395, 84.61029, 82.6452, 78.14883, 72.3955, 69.06921, 61.98898,
    54.39578, 58.4108, 61.42862, 64.58512, 65.65607, 67.33721, 76.59558,
    72.22157, 47.54991,
  51.17789, 53.25573, 55.73647, 58.6202, 61.5108, 67.33811, 77.77771,
    84.44661, 84.37604, 84.24099, 84.28433, 83.92368, 78.99688, 78.51204,
    77.92732, 77.08355, 76.25474, 71.06232, 65.36749, 63.04666, 59.15597,
    57.87282, 61.06615, 63.99031, 65.01192, 64.13481, 67.97414, 73.66646,
    62.05885, 41.40428,
  61.42815, 66.2028, 70.80103, 76.11889, 81.05784, 84.38287, 85.18665,
    84.54116, 79.50111, 77.23097, 72.16588, 66.46625, 62.49603, 61.6632,
    61.2826, 62.00726, 62.5107, 61.0485, 58.7058, 58.22124, 57.80449,
    58.69611, 61.12608, 63.11183, 62.82181, 64.34969, 70.13258, 69.626,
    55.22397, 41.40667,
  72.30913, 75.93955, 78.21555, 80.29396, 83.16326, 82.87718, 71.99157,
    66.34809, 65.45295, 63.64898, 61.88036, 60.81799, 61.50565, 64.97922,
    66.37299, 62.81021, 63.95578, 65.65813, 64.97912, 62.31622, 61.21211,
    64.14841, 67.70206, 67.56936, 66.52112, 72.04071, 74.76137, 63.98231,
    44.17226, 42.12292,
  78.0582, 80.9962, 78.2599, 78.35629, 78.89735, 72.80597, 58.68199,
    62.80766, 63.62761, 66.47786, 69.9159, 73.2169, 72.9138, 71.79723,
    70.1593, 71.63184, 73.03511, 73.07467, 71.48036, 70.8305, 71.24905,
    70.15437, 68.21496, 65.40256, 68.98416, 75.54286, 69.1796, 50.00826,
    41.486, 41.49965,
  76.89912, 77.27448, 77.21466, 76.42458, 79.62151, 73.49484, 67.64393,
    72.81059, 76.75821, 77.53032, 71.64847, 64.22602, 62.92731, 62.90348,
    62.79391, 63.92123, 64.96526, 65.27081, 65.5753, 67.5441, 70.88314,
    68.80827, 63.61407, 63.55066, 68.90417, 66.89814, 51.96567, 41.56252,
    42.16519, 41.37931,
  81.92356, 76.5622, 83.54033, 87.77249, 85.63082, 77.63002, 79.7422,
    73.46622, 67.8996, 67.14399, 62.24808, 59.43119, 60.9833, 60.83903,
    59.09492, 59.53392, 59.20366, 59.55873, 59.93047, 61.69408, 65.63358,
    65.63371, 63.03246, 67.94545, 69.44982, 57.30867, 42.21299, 43.88626,
    42.51877, 41.75393,
  91.04378, 93.83567, 96.46112, 96.84364, 95.35838, 92.13923, 85.19975,
    73.03262, 78.29381, 71.14103, 66.98377, 65.7805, 69.5651, 70.58203,
    65.71798, 57.36049, 58.89685, 59.59711, 59.72851, 61.84147, 65.26769,
    66.05122, 64.14368, 60.08659, 56.78795, 50.61592, 43.49285, 44.76698,
    43.70079, 42.50547,
  94.70483, 96.01143, 95.20902, 92.04279, 89.13462, 87.02444, 85.88327,
    85.59331, 84.30205, 84.3949, 84.55829, 83.74806, 84.26694, 84.67107,
    81.11024, 69.90975, 67.71045, 73.4482, 75.90785, 70.22963, 65.58382,
    60.95399, 55.04274, 49.09195, 45.6702, 44.86332, 43.76788, 43.21242,
    42.96164, 42.34074,
  90.05609, 88.82257, 86.98803, 85.05811, 83.97999, 84.66311, 86.66536,
    86.72177, 85.18053, 84.75146, 84.04797, 81.37337, 81.51431, 83.79688,
    83.58502, 81.92183, 75.99209, 73.60385, 70.91512, 64.86307, 55.81665,
    52.50124, 46.97612, 44.25513, 44.44035, 44.22544, 43.42324, 42.5198,
    41.98236, 41.63787,
  85.79697, 85.60439, 85.61936, 84.42897, 82.98117, 83.38907, 84.16793,
    81.23647, 76.71455, 73.31532, 72.19205, 70.3418, 70.18668, 72.79433,
    70.28813, 68.11249, 66.87933, 61.83107, 57.9921, 53.21214, 48.28278,
    47.21759, 44.36995, 43.81857, 44.18885, 44.06737, 43.19977, 42.47188,
    41.92614, 41.56987,
  76.70007, 75.38911, 74.44904, 73.55098, 72.60549, 71.41068, 71.04163,
    71.12945, 69.05065, 66.63948, 64.21046, 66.31434, 69.03584, 66.13895,
    61.58734, 59.03907, 56.86063, 55.22821, 54.09379, 51.47683, 47.0915,
    47.12412, 44.83062, 43.89276, 44.08965, 44.12149, 43.06978, 42.07333,
    41.76582, 41.55758,
  66.79179, 66.68203, 65.70024, 65.80617, 65.7859, 66.25763, 66.66605,
    67.1252, 66.92444, 65.71877, 67.26171, 68.99692, 67.9564, 65.77196,
    61.33279, 57.79025, 54.76675, 54.27855, 54.49936, 51.67793, 47.0161,
    46.76207, 45.11887, 44.44649, 43.9378, 43.58397, 42.87665, 41.79853,
    41.55096, 41.39516,
  72.61325, 69.17862, 63.26968, 60.06298, 61.14235, 60.98407, 61.28379,
    61.58605, 61.02333, 61.62441, 63.39913, 62.00014, 57.98378, 57.50214,
    56.3421, 57.2379, 61.17158, 64.65709, 64.03072, 59.18966, 52.11843,
    48.14927, 45.70794, 45.01744, 44.15939, 43.45058, 42.78991, 41.84158,
    41.48037, 41.385,
  71.98483, 67.12474, 60.5566, 56.64027, 57.28863, 57.06971, 57.20005,
    57.40115, 58.23351, 60.32257, 60.71839, 57.77901, 57.29087, 56.70165,
    56.18675, 56.96219, 59.74706, 63.01534, 62.88322, 60.06003, 55.35484,
    50.46425, 47.01968, 46.08902, 45.26264, 43.8609, 42.86834, 41.88749,
    41.44831, 41.40691,
  68.80149, 64.35564, 57.97897, 54.54553, 55.07646, 55.10928, 55.60851,
    56.49879, 57.94431, 59.49009, 58.44718, 56.69656, 58.36205, 58.0414,
    56.87331, 56.18108, 56.1933, 56.19068, 55.78038, 54.00701, 52.54441,
    51.47685, 49.30319, 47.81009, 46.36007, 44.36385, 42.86118, 41.94226,
    41.48253, 41.4284,
  67.26418, 63.98175, 57.95566, 55.23969, 55.85658, 55.5798, 56.53536,
    57.48562, 59.25011, 59.49859, 56.62578, 55.0142, 55.72504, 55.14454,
    54.06467, 53.17284, 52.22433, 51.76918, 51.71684, 51.49766, 51.14021,
    50.67081, 50.52197, 49.42097, 47.23827, 44.46437, 42.9507, 42.11541,
    41.56583, 41.43438,
  66.09002, 64.60446, 58.1852, 55.88731, 57.53182, 57.82717, 57.38353,
    56.33814, 56.48146, 55.23251, 52.38401, 52.12016, 52.34122, 52.14915,
    51.34301, 51.33142, 51.21009, 50.47385, 50.20353, 49.90935, 49.53098,
    49.13504, 48.4825, 48.05336, 47.75687, 45.35153, 43.47122, 42.89984,
    42.09294, 41.48603,
  67.66506, 66.97549, 62.40928, 60.72868, 60.98246, 60.0817, 59.93414,
    59.3505, 60.10757, 58.3901, 56.15548, 57.44533, 58.49858, 58.56485,
    57.19961, 56.48773, 55.91604, 54.50611, 52.40795, 51.04737, 50.32941,
    49.68898, 48.6382, 47.89578, 48.04243, 47.55143, 45.6807, 43.66827,
    42.89851, 41.88809,
  69.91912, 67.48084, 61.77184, 59.46681, 59.24212, 58.56631, 59.29915,
    61.70592, 64.89066, 62.9307, 60.13097, 61.80671, 63.00158, 63.19382,
    61.7625, 61.09612, 60.09556, 58.50238, 56.13087, 54.15089, 53.09451,
    51.74005, 49.52812, 48.23006, 48.57151, 48.94704, 48.17418, 45.52011,
    43.99865, 42.79511,
  70.72849, 69.15021, 64.31642, 60.74839, 59.80185, 59.53273, 62.32583,
    66.38115, 67.31195, 63.98621, 63.67868, 64.89758, 65.92703, 65.22114,
    63.19099, 62.44802, 61.53793, 59.87099, 57.59997, 55.78945, 54.88768,
    53.23582, 50.48837, 49.13594, 49.3862, 49.18373, 48.97124, 46.66804,
    43.68482, 42.5762,
  71.68472, 69.87549, 65.67982, 62.81866, 61.97449, 61.21871, 63.90454,
    66.06848, 65.58789, 63.90452, 64.65442, 65.39687, 65.58073, 64.77774,
    63.07992, 62.00257, 61.14971, 59.82916, 58.13205, 57.28531, 57.11742,
    56.64667, 54.97518, 53.34174, 52.62915, 51.63753, 51.13384, 48.86905,
    43.96715, 41.80866,
  72.42838, 71.0248, 67.96002, 66.78777, 67.42176, 66.95271, 67.05145,
    66.41838, 64.59916, 64.38301, 65.04533, 65.73626, 66.28027, 66.30432,
    65.59224, 64.63571, 63.45535, 62.34365, 61.97732, 61.87558, 60.525,
    57.79728, 55.21467, 54.00012, 53.45755, 52.64346, 51.84126, 51.34825,
    48.37223, 43.11839,
  66.32426, 66.40166, 66.53931, 67.03734, 68.88383, 70.71171, 68.63788,
    63.76616, 62.03767, 62.19609, 61.88858, 61.96863, 62.56318, 63.41259,
    63.91425, 63.48561, 62.00805, 60.48226, 58.45563, 56.41178, 54.95567,
    53.45291, 51.77419, 50.64231, 50.45832, 50.08571, 49.11192, 47.60785,
    46.45241, 43.87298,
  61.98402, 62.39767, 62.63297, 62.59215, 64.63095, 68.18472, 68.20406,
    62.70203, 60.04855, 60.88768, 61.22771, 61.63388, 61.11098, 59.79073,
    58.36201, 56.92124, 54.3424, 51.98282, 50.74609, 49.40701, 48.31191,
    48.12563, 47.97237, 47.64206, 47.25031, 46.90675, 45.87857, 44.38685,
    43.15309, 41.7738,
  6.079195, 5.084704, 5.482889, 5.567827, 5.649535, 5.773025, 5.984619,
    6.271905, 6.737524, 7.636083, 9.3976, 11.60629, 13.48307, 17.18169,
    21.45913, 26.31407, 31.92012, 38.55277, 45.53481, 51.55774, 57.63592,
    62.48489, 65.13455, 67.08076, 67.16467, 64.66911, 62.94758, 65.52094,
    59.91935, 57.80554,
  4.537126, 3.775384, 4.077054, 4.572682, 4.844514, 5.064937, 5.432442,
    5.68859, 5.984907, 6.599898, 8.01651, 10.51341, 13.90036, 17.11665,
    21.18041, 26.84916, 33.61473, 40.40876, 46.38574, 52.93746, 58.77071,
    63.88293, 67.63715, 69.97934, 70.83922, 70.19681, 62.59912, 64.03113,
    60.17948, 58.35754,
  7.083001, 6.728895, 7.656177, 8.224352, 9.030512, 9.950092, 10.75697,
    11.4879, 11.99233, 12.35851, 12.86939, 14.11793, 16.26541, 19.32194,
    22.91101, 26.56848, 32.58715, 40.84524, 47.82499, 54.63276, 61.08067,
    66.3243, 69.87792, 71.5443, 71.74464, 71.1288, 70.63566, 65.29254,
    59.15291, 58.3096,
  9.539404, 9.655029, 10.97158, 11.83132, 12.53171, 13.41602, 14.28611,
    15.48039, 16.23476, 16.91637, 18.09422, 19.71553, 21.84942, 24.62212,
    27.86546, 31.49195, 35.25289, 40.2986, 47.85816, 54.65704, 61.35647,
    66.68832, 69.7878, 71.7761, 72.09612, 72.0643, 72.00328, 71.01933,
    66.90773, 58.81811,
  12.07387, 12.4748, 14.12856, 15.08841, 15.60082, 15.77648, 15.92685,
    15.99057, 16.36075, 17.26479, 18.78061, 20.93058, 23.39232, 26.32429,
    29.76955, 33.71566, 38.16674, 43.20842, 49.09748, 55.89474, 61.90907,
    66.27811, 69.62416, 71.46112, 71.9934, 71.99963, 71.77134, 72.54803,
    72.19201, 68.43899,
  11.86923, 12.95229, 15.12085, 16.27253, 16.34457, 16.33982, 16.56299,
    16.71827, 16.75583, 17.23867, 18.55673, 20.70779, 23.77505, 26.89469,
    30.53969, 34.85751, 40.03181, 45.18605, 50.97636, 57.46425, 62.87571,
    64.96239, 70.01882, 71.43045, 71.73362, 71.46722, 71.0402, 71.63682,
    71.62325, 62.45387,
  12.25267, 12.82059, 14.76398, 16.25311, 16.53824, 16.82296, 17.20787,
    17.63765, 17.97986, 18.41606, 19.3649, 20.70264, 18.08275, 22.37901,
    27.47759, 33.83987, 38.90527, 44.90035, 50.78453, 57.53265, 63.2461,
    67.56895, 70.42595, 71.85728, 71.9361, 71.27711, 71.04992, 71.10644,
    70.42134, 56.42839,
  17.00878, 15.85143, 16.35144, 16.4059, 16.5601, 17.01754, 17.39815,
    16.08764, 11.83451, 15.20093, 16.71791, 18.07483, 20.52722, 24.36002,
    28.72232, 33.34568, 38.9976, 45.03965, 51.38191, 57.77468, 63.60898,
    68.0209, 70.76786, 71.86707, 71.75812, 71.5058, 71.59144, 71.11995,
    68.91178, 56.7249,
  19.76535, 17.88355, 17.75214, 17.41932, 17.21632, 17.12795, 16.24468,
    13.46593, 14.01524, 14.82792, 17.16534, 20.23759, 23.54435, 27.00028,
    30.79511, 34.13056, 38.97874, 45.55579, 52.48147, 58.81287, 64.41152,
    68.79974, 71.11507, 71.67956, 71.41664, 71.75967, 71.65646, 70.65641,
    56.91619, 57.27613,
  24.66745, 22.46939, 21.1722, 20.05604, 19.50974, 18.53074, 16.78028,
    17.03722, 17.1056, 17.83957, 19.30736, 22.25184, 25.00441, 27.29074,
    30.08973, 34.82407, 39.81087, 45.53004, 52.03103, 58.97828, 65.25494,
    69.3093, 70.68681, 70.59569, 70.94347, 71.37272, 71.00135, 63.04323,
    56.53479, 56.34947,
  29.68655, 26.64365, 26.67691, 24.30421, 23.20192, 21.40799, 19.87711,
    18.90261, 18.71552, 19.52207, 20.6462, 22.66868, 24.70977, 26.34697,
    29.04769, 33.44958, 38.44963, 44.32697, 51.3343, 57.82932, 64.8005,
    69.09335, 70.44618, 70.65262, 71.00513, 70.70108, 64.48312, 56.9022,
    57.37725, 56.42624,
  30.64736, 27.55497, 30.29502, 30.34595, 29.09068, 25.53153, 22.45446,
    19.63966, 18.56689, 19.30095, 20.71355, 22.76198, 25.85296, 28.43308,
    31.47267, 35.95522, 40.17699, 44.89906, 49.87285, 56.53435, 63.8624,
    68.74892, 70.25513, 71.10628, 71.29662, 70.34711, 57.24923, 60.96272,
    57.91217, 57.03211,
  20.60556, 21.68215, 23.97632, 26.77446, 28.71645, 28.28347, 22.40824,
    17.47779, 20.95364, 20.07306, 21.77855, 23.16585, 25.65402, 28.45139,
    31.84351, 35.3671, 40.38433, 46.00742, 52.19088, 58.48049, 64.09753,
    68.14001, 69.44755, 66.13345, 66.18638, 64.97465, 57.95959, 59.41728,
    58.90956, 57.8117,
  16.91944, 15.55589, 15.23225, 15.94363, 16.47288, 17.27389, 18.25283,
    19.47221, 18.51957, 19.78825, 21.87983, 24.26536, 26.51261, 28.90516,
    32.52017, 36.04698, 39.93221, 46.44336, 53.06892, 59.13619, 63.89782,
    67.48248, 64.36541, 60.41482, 57.64721, 57.9073, 57.3934, 56.98803,
    57.22342, 57.27712,
  17.70189, 11.58867, 14.79599, 15.12505, 16.91916, 17.4455, 17.78265,
    17.94787, 18.46517, 19.93901, 21.93063, 24.37947, 26.97483, 29.8055,
    32.32695, 35.59893, 40.649, 44.96233, 51.94926, 58.65267, 58.75275,
    62.42245, 60.44476, 58.58824, 58.93172, 58.21509, 57.56798, 57.11957,
    56.63401, 56.5697,
  10.03106, 10.96713, 12.69545, 14.55616, 16.36458, 17.68484, 18.32861,
    18.656, 19.27, 21.10933, 23.73745, 26.02604, 28.49217, 30.41275,
    33.13163, 36.56253, 40.34694, 44.65697, 46.85432, 52.35372, 54.18892,
    58.50555, 58.76332, 58.82524, 58.76603, 58.18794, 57.53475, 57.12935,
    56.70414, 56.5723,
  7.388491, 5.687705, 7.187268, 8.662181, 10.44119, 12.72371, 15.30854,
    17.90084, 19.14956, 21.17209, 23.6075, 26.74503, 30.42886, 32.84694,
    35.51986, 38.48139, 41.81227, 45.25121, 49.40538, 53.63664, 54.54656,
    58.54475, 59.07898, 58.8316, 58.75447, 58.38901, 57.52082, 56.72407,
    56.43925, 56.47382,
  10.62259, 7.265922, 6.238048, 6.49048, 7.696902, 8.808593, 10.17222,
    11.69752, 14.15545, 16.938, 21.81049, 25.40737, 28.94599, 33.70608,
    37.71296, 40.83715, 44.26414, 49.55825, 55.95801, 59.85863, 57.69492,
    59.00981, 59.29888, 59.32244, 58.63678, 58.19606, 57.58162, 56.60845,
    56.27942, 56.34077,
  24.41012, 16.3771, 9.211849, 4.039037, 6.047384, 6.241022, 7.246622,
    8.279692, 9.4383, 11.68354, 15.28178, 18.37811, 21.10097, 27.66758,
    35.05213, 40.92738, 46.05028, 52.64693, 59.94148, 65.44914, 66.89382,
    63.03447, 60.76929, 60.7524, 59.42109, 58.64503, 57.87048, 56.76006,
    56.25214, 56.38473,
  23.7872, 16.50566, 9.213462, 4.414557, 5.89332, 6.180421, 7.11188, 8.21699,
    10.03854, 12.99698, 15.52859, 15.97892, 19.23276, 22.40553, 26.54847,
    31.71811, 39.01085, 47.87368, 56.33226, 62.71852, 66.32303, 65.79916,
    62.89457, 62.04887, 60.66394, 59.17442, 58.09992, 56.90306, 56.21634,
    56.36929,
  25.98281, 18.99355, 11.25856, 6.414823, 7.417067, 7.367017, 8.059615,
    8.948971, 10.64557, 12.8099, 14.10602, 15.49681, 19.82075, 23.08858,
    26.52366, 31.23158, 37.27702, 44.41451, 51.68874, 57.58495, 62.32997,
    65.56088, 65.31864, 63.64149, 61.99167, 59.8188, 58.1637, 56.90905,
    56.2289, 56.37622,
  28.03597, 21.99992, 14.73401, 10.81142, 12.27158, 11.83209, 12.35937,
    12.72357, 14.29322, 15.83688, 16.22414, 17.9653, 21.64229, 25.06098,
    28.59214, 33.21703, 38.6859, 44.92091, 51.28682, 56.60776, 60.98398,
    63.74571, 65.35217, 65.38274, 63.74103, 60.75526, 58.77724, 57.45403,
    56.40057, 56.41002,
  28.9209, 24.19882, 17.8096, 14.62094, 17.17228, 18.08874, 18.81243,
    18.81405, 19.73961, 20.68116, 21.70069, 24.89262, 28.3003, 31.68248,
    34.822, 39.01111, 43.89826, 48.69269, 53.84254, 58.29602, 61.8089,
    63.96603, 64.85561, 65.17791, 65.4271, 62.89466, 60.03565, 58.45432,
    57.26794, 56.54815,
  29.00596, 24.53879, 19.53885, 17.4096, 19.36366, 20.06745, 22.1101,
    23.84185, 25.75497, 26.02119, 27.50334, 32.48296, 37.47446, 41.55811,
    44.12498, 47.55426, 51.44489, 55.29817, 59.34201, 63.29686, 66.08574,
    66.99516, 66.53905, 66.09547, 66.3735, 65.94911, 63.39225, 59.83042,
    58.33405, 57.29502,
  28.90198, 23.30606, 17.79852, 14.84251, 16.88056, 17.90092, 19.74044,
    22.40496, 25.05314, 25.80285, 26.63182, 31.53144, 36.88817, 41.38643,
    44.08101, 48.04475, 51.92583, 56.17573, 61.05035, 65.54076, 68.28339,
    68.97536, 67.50925, 66.11047, 66.21653, 65.92381, 65.09262, 61.58311,
    58.91124, 58.02327,
  30.64301, 26.59875, 21.17011, 17.33234, 18.19516, 19.02948, 21.7992,
    24.60316, 25.63005, 26.28115, 29.14732, 33.29365, 38.23064, 41.68699,
    43.88383, 47.53784, 51.67259, 55.93933, 61.13004, 66.00983, 69.23865,
    70.55766, 69.20121, 67.69682, 67.38161, 66.37582, 65.62014, 62.64408,
    58.54396, 57.54967,
  39.13922, 35.54334, 30.74505, 26.884, 27.57758, 27.14155, 29.26772,
    30.65644, 31.13114, 32.22513, 35.62576, 39.60228, 44.00677, 47.10394,
    48.95689, 51.7162, 54.4875, 57.73697, 61.83361, 65.96903, 68.99062,
    70.69582, 70.47243, 69.38705, 69.08624, 68.48541, 68.26231, 65.99734,
    60.31866, 57.13933,
  52.86232, 51.2523, 47.70662, 46.20585, 47.40286, 46.76924, 45.97991,
    45.16989, 44.26367, 45.22637, 46.65073, 49.13208, 52.42034, 54.85394,
    56.24564, 57.74101, 58.63011, 60.21839, 62.8331, 65.96958, 67.24568,
    67.36817, 66.40353, 65.60474, 66.01271, 65.93357, 65.62727, 65.4249,
    63.4531, 58.65847,
  56.17396, 56.90995, 58.63019, 60.82228, 62.5689, 63.98191, 61.84362,
    57.3593, 56.05853, 56.48806, 56.30048, 56.33948, 56.90518, 57.78183,
    58.42163, 58.90338, 58.86366, 58.96203, 59.47991, 60.16568, 61.26563,
    62.3951, 62.48951, 61.85299, 62.03756, 61.9989, 61.42195, 60.12066,
    59.57151, 58.74364,
  60.15104, 60.75882, 61.12058, 61.27599, 62.6976, 65.2655, 65.72029,
    62.09239, 59.83579, 60.62312, 61.11819, 61.54286, 61.54796, 61.02208,
    60.63119, 60.32851, 59.22263, 57.81142, 57.78037, 57.92142, 57.78079,
    58.57727, 59.42895, 59.74529, 59.60799, 59.70429, 59.42175, 58.38549,
    57.42871, 56.62413,
  28.25975, 31.1383, 33.91671, 37.36243, 40.89165, 44.1999, 47.34425,
    50.64644, 54.07582, 57.5743, 61.0845, 64.17819, 66.49613, 68.24759,
    69.42183, 70.07032, 70.31711, 70.33966, 70.23149, 70.01275, 69.53855,
    68.68459, 67.69249, 66.80499, 65.95113, 64.85898, 57.88399, 60.78929,
    56.87307, 54.44855,
  29.2999, 31.60168, 34.16864, 37.21819, 40.64772, 44.19439, 47.86208,
    51.45191, 55.10328, 58.59209, 62.10764, 65.36927, 67.98091, 69.64171,
    70.44868, 70.8101, 70.74013, 70.65424, 70.58144, 70.51885, 70.35483,
    69.97238, 69.29264, 68.49348, 67.71208, 66.19823, 64.52303, 59.035,
    56.26245, 54.76387,
  30.40204, 32.55635, 35.1322, 37.77785, 40.96276, 44.45146, 48.07069,
    51.9916, 55.85697, 59.44501, 62.73301, 65.85525, 68.46828, 70.20654,
    71.1611, 71.3046, 71.02335, 70.74601, 70.45003, 70.22961, 70.29928,
    70.24767, 69.76466, 69.00138, 68.06709, 67.32051, 66.46152, 64.83826,
    56.75601, 54.44905,
  30.91666, 33.43081, 36.11493, 38.8602, 41.69139, 44.72813, 48.13097,
    51.95116, 56.00723, 59.97179, 63.45812, 66.44378, 69.06118, 70.74723,
    71.68734, 72.03436, 71.65787, 71.08017, 70.79853, 70.49146, 70.2735,
    69.71024, 68.41111, 68.10054, 67.37396, 67.38477, 67.54821, 66.79738,
    65.06519, 57.02957,
  31.33844, 33.94344, 37.04937, 40.03785, 42.98819, 45.77457, 48.61595,
    52.18487, 55.71541, 59.63348, 63.34232, 66.64156, 69.57524, 71.44093,
    72.3545, 72.65124, 72.40679, 71.71287, 71.24783, 70.88653, 70.05724,
    68.71836, 67.98223, 67.54842, 67.12296, 66.81283, 66.72636, 67.74185,
    67.35986, 64.87342,
  32.31458, 34.47886, 37.54409, 40.84651, 44.14173, 46.93713, 49.56994,
    53.26608, 56.42935, 59.47453, 62.89093, 66.31953, 69.57361, 71.48541,
    72.66687, 73.11536, 72.79554, 72.29573, 71.45764, 70.88088, 69.86945,
    68.40138, 68.12218, 67.58116, 67.06297, 66.5948, 66.19094, 66.70952,
    66.64592, 59.30519,
  35.25893, 36.22511, 38.5938, 41.18388, 44.31435, 47.41269, 50.22263,
    53.86338, 57.49003, 60.52295, 63.4589, 65.94415, 66.81011, 69.55158,
    70.80405, 71.54498, 71.90305, 71.37154, 70.32665, 69.82269, 69.11842,
    68.4545, 67.96755, 67.65844, 67.1081, 66.57639, 66.43416, 66.4319,
    65.52457, 52.9819,
  40.62026, 40.41019, 41.55497, 43.18766, 45.47782, 48.51511, 51.51434,
    53.26347, 56.05702, 59.32436, 62.22147, 64.8467, 67.30342, 69.40584,
    70.75711, 71.32489, 71.8718, 71.91615, 71.21847, 70.2187, 69.28598,
    68.49374, 67.82988, 67.2447, 66.61689, 66.58516, 66.71792, 66.21408,
    64.59982, 53.2925,
  46.62414, 47.02892, 46.96687, 47.34877, 48.44454, 50.45999, 51.64212,
    54.09074, 57.2953, 60.23508, 62.94044, 65.33563, 67.22528, 69.07141,
    70.54729, 70.83137, 71.43088, 72.12945, 72.22047, 71.29625, 70.20783,
    68.99496, 67.88876, 66.78078, 66.00854, 66.38537, 66.56377, 65.56158,
    53.17177, 53.79718,
  49.89392, 52.80392, 53.76915, 53.54699, 53.20839, 53.37091, 53.52596,
    55.69517, 58.26587, 61.27888, 63.70616, 65.95869, 67.43776, 68.45662,
    69.13941, 70.00963, 70.57512, 71.02895, 71.23402, 71.02339, 70.84845,
    69.40427, 67.72269, 66.26858, 65.83713, 65.88184, 65.55649, 59.95396,
    53.48859, 53.06052,
  48.55877, 51.82944, 56.66417, 58.70746, 58.99649, 57.7578, 57.44886,
    58.16434, 59.60982, 62.57116, 64.67289, 65.98761, 67.25085, 68.1435,
    68.82829, 69.34145, 69.66108, 69.33278, 68.54463, 69.34983, 70.20209,
    69.26511, 67.40067, 66.53728, 66.48577, 65.76776, 63.03954, 54.54,
    54.27589, 53.29439,
  44.76358, 45.02064, 52.68832, 58.54487, 63.51709, 62.65609, 60.29648,
    58.79315, 60.92619, 62.75472, 65.15285, 66.69163, 68.5511, 69.38291,
    69.45863, 69.54041, 69.9418, 70.03384, 69.75146, 69.01571, 69.50605,
    68.98003, 67.05914, 66.32877, 66.27263, 65.38016, 53.49619, 58.8091,
    55.15475, 54.06922,
  38.34374, 41.39992, 44.50206, 50.5949, 57.36528, 62.54966, 61.08012,
    57.7439, 63.64486, 64.48195, 66.95988, 68.4147, 70.07919, 71.13609,
    71.16364, 69.78916, 70.12078, 70.5186, 70.37556, 69.46962, 69.02938,
    68.33852, 67.0176, 62.45472, 61.4128, 62.79198, 54.12944, 55.40303,
    55.80288, 54.83835,
  36.57599, 38.92754, 41.1488, 43.89159, 45.59427, 50.63005, 55.52014,
    60.59755, 62.12494, 65.06702, 67.86115, 70.15493, 71.50663, 72.50031,
    72.4882, 71.25784, 70.42034, 70.59044, 70.90489, 69.60932, 68.175,
    67.0568, 62.60271, 57.72001, 53.93035, 54.13039, 54.16128, 53.27957,
    53.54601, 53.94532,
  34.0185, 31.06915, 39.28722, 43.92576, 47.33387, 50.8223, 53.89614,
    57.45326, 61.76307, 65.13766, 67.63316, 69.71832, 71.58414, 72.94315,
    73.04517, 72.95064, 71.79482, 70.41425, 69.74249, 69.08996, 63.19639,
    63.05017, 58.73861, 55.51627, 55.87414, 54.83931, 54.26732, 53.79091,
    53.26599, 53.2232,
  27.23397, 29.80948, 33.12908, 37.32517, 41.87479, 47.24218, 52.29333,
    55.68075, 59.6425, 63.83132, 67.12296, 69.47404, 71.45733, 73.23766,
    73.83934, 73.64342, 73.41634, 71.99008, 67.99755, 64.20197, 60.28991,
    59.86728, 57.43595, 55.86905, 55.37543, 54.55611, 53.86373, 53.58734,
    53.35522, 53.3002,
  31.06109, 30.02555, 33.27264, 36.49936, 39.8882, 44.1592, 48.47998,
    52.6088, 57.28909, 61.65796, 65.38154, 68.69279, 71.49072, 72.95322,
    73.87105, 74.66576, 75.13517, 74.71663, 73.08637, 69.67681, 62.17759,
    60.36037, 58.19615, 56.24783, 55.57918, 54.89735, 53.88054, 53.28125,
    53.1403, 53.16948,
  41.71606, 37.0901, 36.06362, 37.60854, 41.93748, 45.34342, 49.15937,
    52.88861, 56.37497, 59.35179, 63.96066, 68.44721, 70.55196, 71.83498,
    72.54217, 73.73103, 75.2171, 76.22436, 76.00719, 74.09114, 69.03654,
    62.31846, 59.023, 57.53089, 55.71379, 55.08826, 54.24394, 53.30726,
    53.0709, 53.08327,
  55.06216, 51.14017, 43.62455, 38.7974, 43.79047, 46.66612, 50.58057,
    54.33825, 58.00426, 61.5598, 65.31387, 67.2, 66.75748, 66.94375,
    67.02174, 68.62489, 72.70533, 75.19261, 75.80604, 75.59583, 73.66583,
    67.8396, 61.14704, 59.70122, 57.02699, 55.96014, 54.91928, 53.55595,
    53.05862, 53.1186,
  54.69563, 52.07579, 46.35286, 42.48461, 46.66491, 49.36447, 53.29194,
    57.01904, 60.99427, 64.79106, 67.90175, 69.37029, 71.68953, 70.39788,
    68.76855, 67.48563, 67.89026, 69.91751, 71.14812, 71.88089, 72.37768,
    69.63765, 63.869, 61.20908, 59.01008, 56.92628, 55.36301, 53.7627,
    52.9916, 53.12573,
  56.30251, 53.65474, 49.92946, 46.04409, 50.42886, 52.78791, 56.46486,
    60.30074, 64.52309, 68.10442, 69.64217, 70.40897, 72.96198, 73.73193,
    72.61478, 71.77272, 71.11011, 71.07861, 70.75276, 69.03082, 68.14265,
    67.88744, 65.87636, 62.9381, 60.81494, 58.01306, 55.80698, 53.97099,
    53.00078, 53.09697,
  59.49278, 57.42425, 53.38999, 50.71785, 55.64793, 57.98051, 61.26261,
    64.32576, 68.46587, 72.44518, 74.66432, 76.1051, 77.63292, 78.11969,
    77.29896, 76.00647, 74.42343, 73.15733, 72.07566, 70.50779, 68.79818,
    66.84688, 66.09393, 64.50959, 62.54618, 59.08397, 56.61738, 54.84877,
    53.38582, 53.10875,
  66.29171, 63.56304, 59.92177, 57.07434, 61.49434, 64.07922, 67.25281,
    70.22226, 73.31478, 75.8868, 78.71141, 81.96563, 83.71794, 84.1091,
    83.51936, 82.54956, 81.20377, 78.5127, 76.02357, 73.67911, 71.65807,
    69.05154, 66.67165, 64.91042, 64.44656, 61.44052, 57.80771, 55.96427,
    54.46572, 53.43156,
  75.03867, 72.06921, 67.35085, 64.7085, 67.69237, 68.97884, 71.5118,
    74.3707, 77.41128, 79.55933, 81.82075, 85.20483, 88.37068, 89.46131,
    88.47089, 87.61005, 86.16666, 84.11594, 81.61309, 79.17786, 76.92417,
    73.41155, 69.32557, 66.56683, 65.72989, 64.27243, 61.19103, 57.14033,
    55.44548, 54.30677,
  81.86871, 77.65758, 71.54568, 66.88689, 68.4006, 69.06364, 71.51018,
    74.81963, 77.67677, 79.10735, 80.07762, 83.39151, 86.18074, 87.39568,
    86.42682, 86.03443, 85.24289, 83.72623, 81.49813, 79.35008, 77.5498,
    74.37221, 70.04778, 66.97009, 66.27508, 64.78368, 62.96778, 58.56306,
    55.48366, 54.74195,
  83.85695, 79.30016, 73.94529, 68.4868, 68.39653, 67.73582, 69.88811,
    72.31832, 73.92143, 74.27049, 76.63969, 79.72887, 82.68103, 83.52663,
    82.39078, 82.26839, 81.65523, 79.99022, 78.47699, 77.00136, 75.13026,
    72.88009, 69.36463, 66.80534, 66.43392, 65.2661, 63.86751, 60.29788,
    55.52089, 54.33625,
  80.89805, 77.27874, 72.37242, 67.95364, 68.17749, 66.02798, 66.53858,
    67.54295, 67.61956, 67.32022, 69.33009, 72.39605, 76.31289, 77.78326,
    76.5119, 76.53425, 75.9521, 75.14346, 73.87611, 73.08862, 71.9796,
    70.30663, 67.64789, 65.60562, 65.35938, 64.85466, 64.50405, 62.62813,
    57.77068, 54.38706,
  73.69013, 72.01703, 68.76363, 66.37823, 67.39832, 66.71438, 65.39845,
    64.15614, 62.67332, 62.39485, 62.5577, 63.87925, 66.92023, 68.78892,
    68.51279, 68.43457, 67.78557, 66.92885, 66.66714, 67.3074, 67.04822,
    65.93379, 63.34733, 61.8537, 61.98446, 61.53494, 60.9217, 60.31197,
    59.13728, 55.55974,
  58.84313, 59.75806, 61.155, 62.60634, 63.91406, 65.68464, 64.19201,
    60.3493, 58.77684, 58.96837, 58.44559, 57.90538, 57.85601, 58.66796,
    58.9952, 59.11106, 58.50073, 57.76701, 57.29893, 57.27134, 57.88762,
    58.84312, 59.09536, 58.47538, 58.65327, 58.61287, 57.87516, 56.14766,
    55.35678, 54.96843,
  56.60463, 56.84423, 57.19622, 57.18235, 57.97363, 59.63672, 60.66558,
    58.04068, 56.15922, 56.62775, 56.92908, 56.9894, 56.64801, 56.38548,
    56.37449, 56.2854, 55.59837, 54.39458, 54.09785, 54.05685, 53.8269,
    54.46887, 55.27061, 55.78529, 55.85103, 55.93073, 55.76925, 54.82964,
    53.89044, 53.29514,
  64.05719, 65.57562, 66.52405, 67.34113, 67.75259, 67.99352, 68.12144,
    68.06312, 67.85401, 67.59993, 67.31836, 67.1934, 66.96275, 66.76192,
    66.72974, 66.91033, 67.20398, 67.72486, 68.48135, 69.34831, 70.05236,
    70.60973, 68.1152, 64.41486, 59.5618, 52.28143, 47.47682, 49.80725,
    47.34724, 45.72169,
  63.81318, 65.38905, 66.36266, 67.21651, 67.6777, 67.93895, 68.0542,
    68.12701, 67.97972, 67.67845, 67.42192, 67.23944, 67.16962, 66.96219,
    66.76482, 66.90195, 67.12097, 67.59658, 68.44099, 69.48657, 70.56462,
    71.59765, 72.44273, 72.93354, 72.6734, 66.69067, 50.0707, 47.79194,
    46.74142, 45.81806,
  63.92906, 65.34312, 66.36019, 67.2958, 67.79965, 68.06152, 68.08877,
    68.07458, 67.99142, 67.85544, 67.71117, 67.63759, 67.52445, 67.35418,
    67.33326, 67.28799, 67.39233, 67.74837, 68.31119, 69.21404, 70.41721,
    71.89514, 73.14162, 73.65621, 73.27663, 72.19984, 71.10783, 53.23492,
    46.71902, 45.75897,
  63.99667, 65.32629, 66.2881, 67.25272, 67.92084, 68.31498, 68.34, 68.20231,
    68.07326, 67.84267, 67.82732, 68.09003, 68.09451, 67.8511, 67.81947,
    67.94085, 67.91735, 68.0323, 68.61693, 69.32909, 70.25185, 71.20972,
    65.93406, 70.22222, 70.88211, 72.6429, 72.43421, 71.79198, 58.04351,
    47.78243,
  64.26564, 65.48715, 66.35662, 67.14839, 67.67661, 68.20351, 68.60767,
    68.50793, 68.2589, 67.8959, 67.82409, 68.42514, 68.94024, 68.68796,
    68.65506, 68.72729, 68.73999, 68.73436, 69.07774, 69.71246, 70.12344,
    62.62344, 60.48235, 61.62267, 63.99522, 68.13748, 72.19223, 73.084,
    72.92866, 57.69659,
  64.91111, 65.84605, 66.74396, 67.28353, 67.51773, 67.92355, 68.64531,
    69.02163, 68.89165, 68.46737, 68.27746, 68.64833, 69.21182, 69.18939,
    69.18767, 69.32265, 69.24744, 69.35803, 69.44718, 69.74251, 69.86859,
    59.75912, 63.45622, 63.18418, 63.76546, 64.52531, 66.84099, 72.187,
    72.25838, 50.80264,
  66.70261, 66.66541, 67.34339, 67.76224, 67.92631, 68.23254, 68.73218,
    68.74482, 68.8952, 68.74632, 68.56236, 68.0675, 65.70954, 66.4053,
    66.63296, 67.6608, 68.25158, 68.3391, 66.56158, 66.04483, 63.60779,
    61.38371, 62.86878, 65.06166, 66.42186, 67.33766, 69.4099, 72.26157,
    66.34167, 44.73537,
  70.69606, 69.1548, 68.7726, 68.70139, 68.82464, 69.15775, 69.12426,
    67.67039, 66.73495, 66.77588, 66.13978, 65.57349, 65.61079, 65.80688,
    66.27525, 66.7925, 67.57762, 67.75797, 66.57614, 65.07039, 63.65852,
    63.0631, 63.42044, 64.79567, 66.74652, 70.93479, 72.58764, 70.10295,
    56.83739, 45.00734,
  76.35033, 74.78358, 72.46095, 71.05861, 70.23315, 69.69555, 68.25782,
    67.90852, 67.55865, 67.08472, 66.8292, 66.65646, 65.8579, 66.1058,
    66.67404, 65.95164, 66.95231, 68.61678, 69.79945, 68.94259, 67.54777,
    66.13299, 65.45786, 64.4928, 65.23931, 71.89352, 72.47071, 65.8458,
    44.92738, 45.37936,
  79.69953, 80.85769, 78.98538, 76.37846, 73.89852, 71.54568, 69.0192,
    68.78993, 68.38461, 68.03773, 67.22749, 66.8223, 66.46407, 64.93999,
    63.50062, 63.36322, 63.24372, 63.98082, 65.40267, 67.21136, 68.48769,
    67.83749, 67.18539, 66.32219, 67.90498, 70.24869, 66.50055, 50.2795,
    44.9856, 44.93375,
  77.83519, 80.40896, 83.47153, 82.59757, 80.31164, 75.52242, 72.2697,
    70.32861, 69.23824, 69.34766, 68.05345, 66.75401, 66.3939, 66.29318,
    63.47201, 63.05336, 61.29056, 59.81517, 59.86522, 61.21844, 64.05385,
    64.64075, 64.85492, 70.24342, 72.1897, 72.01492, 53.32513, 45.79537,
    45.88344, 45.08966,
  73.47933, 73.5979, 79.15325, 83.04111, 83.9558, 80.21503, 75.25059,
    71.49593, 70.27012, 69.66843, 68.80019, 67.78088, 67.61333, 67.33332,
    66.80303, 66.78946, 66.94602, 64.07837, 60.92817, 59.53073, 61.52678,
    61.90367, 60.14389, 63.68159, 70.86668, 67.69944, 45.37647, 50.14886,
    46.68618, 45.74057,
  67.28276, 69.09712, 70.76483, 74.06316, 77.42214, 78.90844, 74.27885,
    70.37617, 72.49088, 71.09854, 70.44358, 69.36237, 69.12755, 68.84196,
    68.12694, 66.89995, 67.48631, 68.4301, 69.16808, 63.81734, 62.99585,
    63.30248, 59.76797, 53.72881, 52.20167, 53.48565, 45.81536, 47.27819,
    47.45862, 46.45723,
  68.13448, 68.66946, 68.03871, 65.47436, 64.80418, 68.53442, 70.65475,
    72.05302, 70.40675, 71.0591, 71.14722, 70.63619, 70.26642, 69.90496,
    69.02692, 67.79678, 67.27823, 68.09956, 69.28177, 69.5826, 64.57446,
    60.74487, 52.98219, 48.79622, 45.38942, 45.60439, 45.7042, 45.07518,
    45.38755, 45.69942,
  68.65114, 66.6269, 69.71259, 69.49886, 69.33916, 69.29398, 69.66595,
    69.80721, 69.79901, 69.60983, 69.78788, 69.90167, 70.2354, 70.22961,
    69.50398, 68.92324, 68.00879, 67.45784, 64.96854, 61.77999, 54.6488,
    53.92877, 50.0279, 46.75833, 47.06088, 46.2884, 45.8724, 45.42334,
    45.05773, 45.07237,
  64.29613, 66.85475, 67.64166, 68.4054, 68.18206, 69.14162, 70.02174,
    69.96133, 69.41995, 69.00872, 69.20204, 69.68754, 70.31921, 70.93128,
    70.50232, 69.78331, 69.40137, 66.38165, 59.61289, 56.54974, 53.22917,
    51.46292, 48.63403, 47.03848, 46.58649, 46.0069, 45.53996, 45.31985,
    45.13186, 45.11479,
  68.00694, 67.70493, 68.58834, 69.27771, 68.96922, 68.31283, 68.42422,
    69.30811, 69.17092, 68.3593, 68.69819, 69.38644, 70.4653, 70.84299,
    70.9434, 71.19236, 71.32814, 71.07603, 65.89419, 60.73334, 54.40294,
    52.4226, 49.79827, 47.53536, 46.89817, 46.31008, 45.5141, 45.04333,
    44.99432, 45.02172,
  77.11245, 73.47125, 70.70399, 70.43536, 71.17022, 70.74638, 70.55779,
    70.00904, 69.96732, 68.36735, 68.27311, 69.09109, 69.79097, 69.70637,
    69.80745, 70.67938, 71.76833, 72.76881, 73.12537, 68.7317, 60.02929,
    53.91186, 50.86721, 48.97044, 47.35576, 46.70135, 45.84649, 45.0764,
    44.93505, 44.95882,
  87.6515, 82.9613, 75.86871, 70.09002, 72.56361, 72.17928, 71.93094,
    71.3748, 70.62865, 70.43129, 70.27415, 68.84969, 66.30758, 63.86424,
    61.88329, 62.67695, 66.20562, 70.544, 72.28318, 72.42896, 66.93835,
    58.42516, 52.47598, 51.03589, 48.61718, 47.63829, 46.58037, 45.32884,
    44.92218, 44.95811,
  85.99686, 82.29588, 75.66426, 70.82028, 73.09334, 73.4069, 73.53206,
    72.89687, 72.53802, 72.62025, 72.17918, 71.20983, 70.87428, 67.55376,
    63.93003, 61.98005, 61.5654, 62.69492, 63.179, 63.33627, 62.91003,
    59.56336, 54.54956, 52.18497, 50.19631, 48.43233, 46.99663, 45.51848,
    44.85007, 44.96318,
  84.96159, 81.68314, 75.41185, 70.65264, 72.89389, 73.48612, 74.34461,
    74.56335, 74.99243, 74.59801, 72.85579, 70.91358, 71.01857, 70.35098,
    68.24785, 66.80375, 65.67067, 64.71571, 63.29899, 60.74176, 58.91415,
    57.96318, 55.97505, 53.10761, 51.41159, 49.22358, 47.27394, 45.60785,
    44.80463, 44.96541,
  82.11113, 80.07086, 73.79193, 69.8768, 72.3744, 73.02783, 74.37972,
    75.20684, 76.67458, 77.66464, 76.51739, 74.56311, 73.42473, 72.60096,
    71.35738, 69.89256, 68.38322, 66.9709, 65.21941, 62.69402, 59.91935,
    57.24519, 56.74852, 53.94228, 52.55617, 50.11438, 48.00016, 46.2546,
    45.05212, 44.92905,
  80.20744, 77.42428, 72.49799, 68.48028, 71.4139, 72.85248, 74.48913,
    75.3755, 77.03834, 78.43186, 79.07298, 79.3746, 79.18379, 78.73882,
    77.43385, 75.8466, 73.71587, 71.17701, 68.85195, 65.99056, 62.99136,
    59.7005, 57.51553, 54.98539, 54.099, 51.92178, 49.06011, 47.25337,
    45.88185, 45.13148,
  79.2143, 76.21664, 71.03931, 67.93626, 69.81675, 70.97198, 72.78551,
    74.68066, 76.73946, 78.02208, 79.40163, 81.16489, 83.07174, 83.78593,
    82.71934, 81.99816, 80.53583, 76.95477, 74.02384, 71.25203, 68.13747,
    64.34643, 60.02982, 56.98007, 55.98075, 54.51433, 51.82361, 48.41498,
    46.76942, 45.86053,
  79.58873, 75.50586, 68.91884, 64.29122, 65.17519, 65.62185, 68.04373,
    71.38306, 75.14512, 75.79173, 76.53299, 79.0899, 82.00317, 83.19917,
    81.24755, 80.73232, 78.66663, 76.56647, 73.95518, 71.74341, 68.70798,
    65.21534, 60.67899, 57.56839, 56.6156, 55.19708, 53.58519, 49.55138,
    46.97831, 46.32504,
  80.50558, 74.99927, 67.65575, 62.34161, 62.16704, 61.48374, 63.28796,
    66.18962, 68.73086, 69.5149, 71.69813, 74.41749, 77.14405, 78.00114,
    76.0513, 75.09028, 74.5307, 72.29153, 70.58778, 69.08675, 66.80136,
    64.04942, 60.26539, 57.52391, 56.93046, 55.71049, 54.37003, 50.94566,
    47.01118, 45.95901,
  75.53421, 71.82092, 64.73961, 60.28936, 60.48693, 58.62043, 58.88722,
    59.99198, 60.93992, 61.24208, 63.4898, 66.39404, 69.84737, 71.07216,
    69.52005, 68.95802, 68.49049, 67.24686, 66.03181, 64.96086, 63.56049,
    61.36212, 58.58435, 56.52489, 56.16698, 55.40112, 54.84034, 52.51736,
    48.55942, 46.01157,
  64.99968, 64.24541, 59.99754, 57.24415, 58.65247, 58.21154, 56.68566,
    55.78819, 54.84931, 54.75632, 55.17998, 56.83293, 59.72132, 61.48684,
    61.127, 60.91825, 59.94083, 58.93306, 58.65806, 59.0616, 58.45543,
    57.10405, 54.6288, 53.36859, 53.36086, 52.94619, 52.25029, 51.00886,
    49.60463, 46.88537,
  50.17297, 51.29774, 52.35346, 53.27943, 54.36688, 55.97106, 54.73961,
    51.6705, 50.42222, 50.51141, 50.14363, 49.8278, 49.88258, 50.53843,
    50.71928, 50.76925, 50.32773, 49.62988, 49.15316, 49.3353, 49.80215,
    50.5575, 50.83422, 50.143, 50.25107, 50.23748, 49.48029, 47.81209,
    46.94001, 46.34587,
  47.84945, 48.12967, 48.44093, 48.43685, 48.9869, 50.38814, 51.1996,
    49.25552, 47.82594, 48.20406, 48.37764, 48.42096, 48.23867, 47.95004,
    47.92696, 47.88695, 47.18649, 46.14908, 45.95592, 45.918, 45.80661,
    46.40911, 47.3139, 47.68195, 47.487, 47.55286, 47.44872, 46.49673,
    45.64498, 45.15643,
  62.65215, 62.75131, 62.90867, 63.11456, 62.92078, 62.422, 61.58665,
    60.56467, 59.54833, 58.79986, 58.53555, 58.6528, 58.73188, 59.68162,
    61.19542, 62.80492, 64.32692, 65.39845, 64.55025, 62.94317, 61.501,
    60.3186, 58.47985, 56.70934, 54.41076, 50.58453, 47.93901, 49.54295,
    47.41592, 46.11072,
  64.62506, 64.65356, 64.44959, 64.72597, 64.74685, 64.79635, 64.73663,
    64.15369, 63.10828, 61.81118, 60.63057, 59.79628, 59.24486, 58.85034,
    59.17965, 60.63592, 62.84055, 65.89284, 65.33228, 63.98763, 62.7442,
    61.75154, 61.0387, 60.75669, 60.36136, 58.86372, 48.87992, 47.80682,
    47.12547, 46.16028,
  65.52676, 66.11603, 65.98046, 65.71066, 65.27906, 65.15694, 65.31804,
    65.67551, 65.85396, 65.57143, 64.73949, 63.67211, 62.55661, 61.62425,
    60.67474, 59.45031, 59.25749, 60.52731, 63.31555, 64.00163, 63.2351,
    62.61722, 62.15469, 61.73124, 60.97157, 59.95487, 59.21542, 50.89946,
    46.63369, 46.23708,
  65.9384, 66.87963, 67.78492, 68.36607, 68.20609, 67.60091, 66.85547,
    66.44861, 66.93995, 67.69892, 68.60085, 69.28571, 68.4304, 66.90561,
    66.20563, 65.1534, 63.33692, 61.63541, 61.81638, 63.65069, 63.16796,
    62.25799, 61.12244, 61.04801, 60.62722, 60.8042, 60.26295, 59.74613,
    55.10163, 47.61484,
  66.75043, 66.63139, 67.65966, 68.83664, 69.48357, 69.97379, 70.42869,
    69.46903, 68.14323, 67.78398, 69.48582, 70.66271, 71.13863, 70.47605,
    69.75255, 69.1102, 68.05804, 66.64319, 65.15102, 63.46461, 62.29963,
    59.2293, 57.38447, 59.48465, 60.55021, 60.24625, 60.32571, 61.18204,
    61.14135, 56.70742,
  68.18339, 68.10668, 67.85587, 68.24469, 69.09708, 70.09893, 71.07246,
    71.61534, 71.50248, 71.16833, 71.08187, 71.51556, 71.79153, 70.77367,
    70.01897, 69.19772, 67.69179, 67.00549, 66.30751, 64.67207, 63.02486,
    56.55495, 60.16539, 59.86222, 59.97353, 59.76038, 59.92193, 60.24252,
    60.38958, 51.75102,
  68.67222, 68.7663, 68.9352, 69.0275, 69.31154, 70.15775, 71.22804,
    71.93478, 72.30793, 72.07868, 71.95023, 71.48566, 60.24274, 60.10888,
    59.50089, 59.90218, 61.92918, 61.61232, 59.81794, 60.22866, 59.003,
    58.52585, 60.70127, 60.85728, 60.67541, 60.52288, 60.57129, 60.3725,
    59.45911, 45.20868,
  70.22478, 69.59381, 69.5211, 69.50803, 69.74894, 70.46677, 71.01999,
    62.93048, 56.49005, 58.7215, 58.87334, 58.78301, 59.10992, 59.65346,
    60.18779, 60.40881, 60.27018, 59.7051, 58.57065, 57.71106, 57.66312,
    58.38222, 60.12564, 60.58257, 60.55966, 60.87671, 60.96755, 60.26542,
    57.38995, 45.39144,
  73.89252, 72.48904, 71.34911, 70.80731, 70.69007, 70.73374, 66.3409,
    62.12901, 60.12863, 58.03042, 57.50719, 57.67326, 57.94193, 59.56008,
    61.19143, 61.09052, 62.12288, 63.43018, 63.85107, 62.5976, 61.39159,
    60.9375, 60.62788, 59.99406, 60.05478, 60.86941, 61.13706, 59.96206,
    45.47223, 45.87176,
  78.94572, 77.99277, 75.97363, 74.21629, 73.08932, 71.68002, 70.05701,
    70.33745, 67.45122, 63.71267, 59.54197, 57.81937, 56.72017, 55.73637,
    55.69973, 56.895, 58.43447, 60.19068, 61.94269, 63.4096, 64.22868,
    62.32982, 60.65815, 59.65795, 59.76508, 60.073, 59.95976, 50.55954,
    45.40496, 45.45312,
  82.0873, 82.05128, 82.64094, 80.13886, 78.11032, 74.65778, 72.4769,
    71.19127, 70.62164, 70.81401, 67.86664, 60.72319, 57.80637, 55.21918,
    53.56875, 53.78073, 53.73247, 54.38749, 55.854, 58.04174, 61.69766,
    62.41299, 60.55943, 60.13526, 60.66411, 60.32532, 52.41363, 45.7767,
    46.24102, 45.5279,
  81.1728, 80.55717, 83.94939, 85.14584, 83.66877, 79.63102, 75.57217,
    72.19324, 70.74892, 70.65094, 69.72866, 68.66412, 67.88542, 65.64757,
    60.20636, 57.09071, 56.95325, 55.80223, 54.85494, 55.22392, 58.11163,
    59.37593, 58.4064, 59.91494, 60.14908, 59.68544, 45.95163, 49.81377,
    46.91014, 46.03276,
  72.36443, 74.49107, 76.59218, 79.31811, 81.33718, 81.15841, 75.54913,
    71.08606, 73.03044, 71.58555, 70.80352, 69.8174, 69.45143, 68.98842,
    67.83051, 61.38154, 63.56522, 64.21997, 62.4981, 58.35034, 58.92405,
    60.17947, 57.98393, 53.09816, 52.16841, 53.11209, 46.13874, 47.81207,
    47.71134, 46.70231,
  70.63275, 68.03629, 64.4379, 62.74233, 63.36861, 70.12324, 72.77217,
    73.35526, 71.23315, 71.71637, 71.4022, 70.19667, 69.72643, 69.48254,
    68.16916, 66.65453, 65.72247, 64.93248, 64.2454, 62.61758, 60.66667,
    57.46924, 50.71054, 47.77974, 45.67894, 45.98599, 45.9777, 45.55952,
    45.96547, 46.1345,
  69.3249, 65.0283, 65.85971, 64.40983, 63.69492, 63.65141, 64.79368,
    64.81891, 64.53593, 64.05, 64.04312, 63.3382, 65.39016, 66.85872,
    68.24456, 67.9355, 66.51079, 62.15469, 60.03457, 56.91126, 50.8367,
    51.48207, 49.1669, 46.21679, 46.94404, 46.64727, 46.1625, 45.70953,
    45.49866, 45.53996,
  61.2931, 62.87236, 63.22289, 63.43817, 63.27469, 64.14493, 65.285,
    65.99877, 65.04723, 63.92025, 63.96213, 63.89181, 64.25544, 65.27661,
    62.35246, 60.83048, 61.0606, 56.39853, 52.41468, 51.01796, 49.38819,
    48.92183, 47.21542, 46.39844, 46.54211, 46.48979, 46.04049, 45.73404,
    45.60349, 45.60987,
  62.54668, 61.3001, 61.04905, 60.89165, 60.3651, 59.99443, 60.77355,
    62.59684, 63.42788, 63.25862, 63.6212, 66.25881, 69.79187, 70.09544,
    66.24303, 64.26828, 62.00132, 59.49472, 56.03054, 53.03983, 49.56597,
    49.2148, 47.71518, 46.73954, 46.82238, 46.65955, 45.9396, 45.50887,
    45.51326, 45.55097,
  69.32375, 65.50599, 62.32604, 61.17259, 60.62903, 59.76335, 59.59063,
    59.81806, 60.18171, 59.52944, 60.70809, 62.50069, 64.71779, 66.61765,
    65.91192, 66.75315, 67.42897, 66.363, 64.10091, 59.64529, 53.61412,
    50.21878, 48.59514, 47.83318, 47.32338, 46.96885, 46.1878, 45.52571,
    45.48003, 45.50793,
  84.23483, 76.79324, 67.26648, 61.30005, 62.07488, 60.86456, 60.43421,
    59.98321, 58.89235, 58.35461, 58.16963, 57.23857, 55.62791, 55.20156,
    55.34533, 57.39189, 61.40965, 65.6956, 66.81659, 65.57556, 60.36985,
    53.99187, 50.26957, 49.66647, 48.41279, 47.86803, 46.9094, 45.77843,
    45.51061, 45.51447,
  83.51942, 77.324, 68.80565, 63.54567, 64.12897, 63.28624, 62.80773,
    61.96037, 61.36008, 61.02385, 60.43174, 59.2298, 58.44593, 55.21283,
    52.94138, 52.27705, 53.45375, 56.02055, 57.8033, 58.34418, 58.0136,
    55.46519, 51.91051, 50.87719, 49.7079, 48.50988, 47.28248, 45.99697,
    45.45012, 45.53802,
  83.40521, 78.82336, 69.94002, 65.51226, 66.27452, 65.72568, 65.53989,
    65.02, 64.41216, 63.22327, 61.42709, 60.01667, 60.14196, 58.90725,
    56.64914, 55.84723, 55.69672, 55.93731, 55.69492, 54.30909, 54.00602,
    54.23216, 53.25828, 51.66727, 50.70908, 48.92992, 47.33479, 45.94986,
    45.45251, 45.54865,
  80.11172, 78.17056, 69.6113, 66.1132, 67.72634, 67.68076, 68.13512,
    68.30607, 68.6858, 68.11824, 66.06962, 63.93596, 62.7296, 61.55101,
    60.1567, 59.04654, 58.27008, 57.90888, 57.13834, 55.4493, 53.49923,
    52.69512, 54.09526, 52.33069, 51.79214, 49.76794, 47.87035, 46.31846,
    45.54282, 45.49104,
  77.57304, 75.22075, 67.74786, 64.95748, 67.17532, 68.09577, 69.02129,
    69.77944, 71.33366, 71.92458, 71.34483, 70.9292, 70.02141, 68.84657,
    66.99987, 65.36014, 63.81061, 62.51325, 61.2169, 59.00866, 56.41949,
    54.49905, 54.7213, 53.46552, 53.53136, 51.59904, 49.08077, 47.16792,
    46.14262, 45.62898,
  74.8056, 71.66659, 65.54027, 63.44667, 65.09113, 65.75666, 67.4227,
    69.70364, 72.72424, 73.90971, 74.10122, 76.02879, 77.87266, 77.94479,
    75.7967, 74.08835, 71.63903, 68.76028, 66.91648, 64.72347, 62.23409,
    59.4959, 56.71314, 55.44156, 55.26428, 54.23074, 51.81003, 48.53915,
    46.96305, 46.11335,
  73.82394, 68.62894, 62.11299, 58.92454, 59.87245, 60.50858, 63.04661,
    67.07655, 71.37509, 71.48741, 71.12011, 73.42232, 76.1096, 76.93446,
    74.86834, 73.56999, 71.47433, 68.77786, 67.53201, 66.28459, 63.63745,
    60.90553, 57.84488, 55.8726, 55.77659, 54.7575, 53.23552, 49.7271,
    47.23718, 46.5257,
  73.02576, 68.12268, 61.87255, 57.48537, 57.51594, 57.2053, 59.55135,
    63.57348, 67.00314, 67.35386, 68.66393, 70.76624, 73.63377, 74.49747,
    72.82467, 71.41652, 69.80647, 67.41058, 66.15893, 65.3831, 63.40486,
    61.02825, 58.4016, 56.83094, 56.26656, 55.06055, 53.86254, 50.67641,
    47.13133, 46.27364,
  70.95728, 67.18443, 61.33135, 57.45129, 57.49546, 55.96916, 56.6892,
    58.61024, 60.69308, 61.23417, 63.16356, 65.77947, 68.84642, 70.23321,
    69.44621, 68.64102, 67.29486, 65.34103, 64.15853, 63.45749, 61.91478,
    59.88494, 57.79724, 56.3717, 56.24977, 55.26032, 54.90857, 52.55445,
    48.31557, 46.22779,
  64.79706, 63.29787, 59.38373, 56.93056, 58.09312, 57.30948, 56.02422,
    55.73209, 55.15412, 55.29645, 55.91872, 57.84575, 60.64748, 62.30985,
    62.23801, 61.91434, 60.83595, 59.72615, 59.58493, 59.77403, 59.09937,
    57.28857, 54.81284, 53.56824, 53.53011, 53.17122, 52.5743, 51.5373,
    49.79909, 47.01175,
  51.39245, 52.42426, 53.17363, 53.96511, 55.42186, 57.04533, 55.33403,
    51.98829, 51.00397, 51.24789, 50.82293, 50.64982, 50.78392, 51.36218,
    51.31071, 51.17762, 50.94915, 50.59711, 50.13096, 50.42789, 50.90324,
    51.46922, 51.26052, 50.53537, 50.56994, 50.45201, 49.71358, 48.18925,
    47.48851, 46.78952,
  48.52858, 48.7132, 49.12637, 49.2751, 50.15813, 52.00779, 52.61207,
    49.99766, 48.5436, 49.07889, 49.4751, 49.43192, 49.17606, 48.79279,
    48.65339, 48.43782, 47.59953, 46.77799, 46.64117, 46.66528, 46.65369,
    47.22066, 47.94727, 48.17965, 48.14293, 48.22962, 47.90227, 46.94772,
    46.23466, 45.70568,
  56.50787, 56.46486, 56.19626, 56.01447, 55.62376, 55.38121, 55.31388,
    55.34487, 55.59086, 56.15942, 57.11777, 57.85803, 57.81802, 57.61562,
    57.07001, 56.23033, 55.27917, 54.2907, 53.26638, 52.06463, 50.00422,
    47.72799, 46.65875, 46.6182, 46.07751, 43.25564, 41.26736, 42.65178,
    39.13979, 37.61035,
  60.29464, 60.53313, 60.10576, 60.03646, 59.52113, 59.02453, 58.64917,
    58.17247, 57.69686, 57.3971, 57.54964, 58.28342, 58.82197, 58.36998,
    57.77495, 57.12756, 56.32007, 55.48163, 54.58548, 53.67444, 52.88462,
    52.22555, 51.84641, 52.02047, 52.09725, 50.84871, 39.58685, 41.16089,
    38.99596, 37.8515,
  61.51235, 62.10734, 62.13811, 62.15421, 62.09445, 62.19767, 61.82441,
    61.34935, 60.7707, 60.14637, 59.58689, 59.12593, 58.28011, 57.85155,
    57.68231, 56.84597, 56.1204, 55.60456, 55.06507, 54.42293, 54.09787,
    53.928, 53.74392, 53.51303, 52.88588, 51.47804, 50.27794, 41.81549,
    38.47924, 38.00595,
  63.20919, 64.19871, 64.53186, 64.14762, 63.48694, 62.87831, 62.37501,
    61.74636, 61.05676, 60.29445, 59.85935, 59.87569, 59.57877, 58.74126,
    58.16108, 57.42062, 56.29451, 55.5318, 55.19559, 54.79918, 54.36216,
    53.67297, 53.36773, 53.6947, 53.13079, 52.23378, 51.46252, 50.72364,
    43.82527, 38.71369,
  63.80568, 65.37959, 64.93491, 64.45901, 63.77547, 63.302, 62.95282,
    62.12585, 61.12609, 60.05147, 59.71125, 60.35334, 60.67273, 60.03014,
    59.42745, 58.94007, 57.70795, 56.07768, 55.27604, 54.96588, 53.8849,
    52.46167, 52.32905, 52.85398, 53.02031, 52.59224, 52.41006, 52.92302,
    52.4332, 46.92116,
  62.5751, 65.12746, 65.09216, 64.53535, 63.7715, 63.697, 64.17154, 63.62029,
    62.5704, 61.49027, 60.96333, 61.24852, 61.50005, 60.85087, 60.77634,
    60.30795, 58.70767, 57.25445, 55.37988, 54.59077, 53.41076, 49.63597,
    52.27492, 52.42517, 52.51742, 52.64583, 52.86387, 53.56438, 52.51297,
    41.31435,
  61.98824, 63.67424, 64.82528, 64.37728, 63.84752, 64.03698, 64.81681,
    64.76714, 64.02169, 62.87125, 61.93792, 60.71798, 58.73073, 58.9577,
    58.5512, 57.84842, 56.97738, 55.75426, 54.55436, 53.90407, 52.96925,
    52.37644, 52.38061, 52.62927, 52.44378, 52.25439, 52.83116, 52.89504,
    51.09159, 36.76798,
  64.44063, 64.25353, 64.10063, 63.89417, 63.59703, 63.83781, 64.18106,
    63.05376, 61.07777, 61.59792, 60.92633, 60.29451, 59.41636, 58.94262,
    58.46784, 58.01542, 57.23293, 56.28953, 55.24442, 53.98147, 53.07625,
    52.68664, 52.62509, 52.59845, 52.32341, 52.56764, 53.17601, 52.57507,
    48.45927, 36.98124,
  65.2418, 64.59831, 63.89313, 63.40291, 62.87139, 62.44725, 59.68497,
    58.69929, 59.85517, 60.04911, 60.67738, 60.3188, 59.99358, 59.99759,
    59.75499, 58.76633, 58.3568, 57.91852, 56.96465, 55.31985, 53.91637,
    53.17458, 52.83902, 52.30585, 52.19729, 52.87504, 52.70139, 51.38862,
    37.33273, 37.51952,
  67.89814, 67.09406, 65.7371, 64.71455, 63.77653, 62.19017, 58.95195,
    60.40654, 59.16572, 57.85287, 56.97296, 57.78118, 57.76395, 57.44993,
    57.27288, 57.63244, 57.64157, 57.48371, 56.94783, 56.28573, 55.40434,
    53.65467, 52.25321, 51.43571, 52.12975, 52.81059, 51.77314, 42.62267,
    36.9939, 36.90158,
  72.26738, 70.82487, 71.1342, 68.4668, 67.42882, 64.00517, 61.83841,
    60.31474, 59.47268, 58.88857, 56.64522, 51.92018, 51.55573, 50.6031,
    49.91772, 50.30777, 51.10558, 52.08103, 53.80714, 54.85731, 55.16764,
    53.78991, 51.92495, 51.57322, 52.04745, 51.68724, 44.55149, 37.35293,
    37.94278, 36.9995,
  77.18819, 75.40501, 76.52306, 76.17547, 72.85305, 68.6205, 64.82895,
    61.43907, 59.53233, 59.03619, 57.77929, 56.47586, 55.81601, 56.09036,
    55.02008, 51.84532, 51.48388, 50.67948, 50.33469, 51.46388, 54.17579,
    53.53544, 51.82516, 51.98294, 52.12145, 50.9116, 37.87248, 41.53398,
    38.49321, 37.5367,
  69.11223, 71.14444, 72.57629, 73.84315, 74.01084, 71.93144, 65.04453,
    60.54107, 61.74221, 59.88286, 58.80712, 57.76581, 57.36786, 57.28906,
    56.87178, 55.14742, 54.97916, 54.66108, 54.16732, 52.94106, 53.67357,
    53.19821, 51.77708, 47.64705, 47.12395, 45.08674, 38.28401, 39.88976,
    39.51167, 38.23294,
  64.40328, 64.20119, 64.06857, 62.54066, 62.10254, 62.49851, 63.00889,
    62.61482, 59.98775, 59.94534, 59.30291, 57.73892, 57.41357, 57.32488,
    56.39994, 55.73101, 55.50948, 55.12282, 54.9558, 53.85006, 53.197,
    52.31866, 46.71855, 40.41396, 37.5019, 37.98035, 37.65027, 37.37966,
    37.77539, 37.72333,
  67.23184, 63.60398, 64.12045, 62.60996, 61.88028, 61.78919, 62.78072,
    62.25115, 60.19417, 58.98397, 58.27313, 57.7379, 57.82713, 57.14989,
    56.82769, 56.94061, 55.45893, 55.40427, 54.90908, 53.75253, 48.00452,
    45.22865, 40.54171, 38.56752, 38.9946, 38.46504, 37.85947, 37.46498,
    37.15496, 37.06997,
  59.58015, 62.55445, 63.58881, 64.41252, 64.87157, 64.84796, 64.6114,
    63.69487, 62.00047, 60.00415, 59.04206, 58.1963, 57.7589, 57.95373,
    56.87403, 55.68643, 55.60409, 51.89918, 48.19458, 45.50118, 42.19224,
    41.39966, 39.22646, 38.43927, 38.62125, 38.43928, 37.84249, 37.4857,
    37.27526, 37.13277,
  56.2938, 56.40191, 57.40183, 58.6162, 59.73437, 60.93667, 62.84457,
    64.21799, 63.42757, 61.92777, 60.47751, 60.26151, 60.57984, 59.84853,
    58.1776, 57.59641, 55.20735, 53.23742, 50.68121, 47.30149, 42.95596,
    41.94903, 39.73046, 38.71216, 38.79162, 38.61718, 37.69235, 37.09903,
    37.08169, 37.08607,
  60.86748, 58.34411, 56.07725, 55.83028, 56.38479, 57.18317, 58.7047,
    60.79799, 62.42522, 62.86335, 62.33204, 62.00079, 61.52098, 60.70818,
    59.76254, 59.81719, 60.2048, 60.06903, 58.50057, 53.34694, 46.24702,
    42.94228, 40.75867, 39.7452, 39.09384, 38.59296, 37.83514, 37.00798,
    36.97008, 36.98791,
  76.31723, 69.17931, 59.48137, 53.92061, 55.01162, 54.61293, 55.30908,
    56.07379, 56.31361, 57.18157, 58.47155, 58.16388, 56.48521, 56.42643,
    56.20652, 58.0839, 60.28839, 61.56398, 60.79371, 58.85663, 53.52668,
    46.6318, 42.86546, 41.70692, 40.37066, 39.37204, 38.31587, 37.2276,
    36.94294, 36.99871,
  76.86498, 70.37727, 61.27755, 55.98407, 56.50549, 56.09123, 56.18644,
    56.29324, 56.67717, 57.53128, 57.38413, 55.75467, 55.38345, 52.88252,
    50.66075, 50.1019, 51.649, 54.60658, 55.84366, 55.04258, 52.67236,
    48.58769, 44.72998, 43.10926, 41.70299, 40.05109, 38.71455, 37.39492,
    36.91401, 36.99876,
  78.94009, 73.68622, 64.701, 59.70543, 59.90987, 59.14359, 58.96874,
    58.72002, 58.72126, 58.591, 57.15322, 55.82284, 56.47298, 55.53118,
    53.68099, 52.84367, 52.65039, 52.67191, 52.18669, 49.97417, 48.64568,
    47.81226, 45.86934, 44.23157, 42.67901, 40.56062, 38.8397, 37.45504,
    36.92308, 37.00103,
  79.16481, 76.71338, 68.63325, 64.53342, 65.20434, 64.30766, 64.17876,
    63.72387, 63.731, 62.90065, 60.7335, 59.00584, 58.28106, 57.21563,
    55.88258, 54.95411, 54.0246, 53.4226, 52.67462, 51.26668, 49.64916,
    47.32035, 45.90639, 45.01551, 43.68902, 41.26246, 39.28992, 38.04559,
    37.08461, 36.95896,
  78.77347, 77.38898, 70.18906, 67.26262, 68.8531, 69.16424, 69.34412,
    69.15894, 69.85079, 69.38973, 67.86918, 67.5627, 66.40846, 64.57045,
    62.41273, 60.70189, 58.70051, 56.37904, 54.58259, 52.55167, 50.60736,
    48.24789, 46.00111, 45.46824, 45.53533, 43.24771, 40.42078, 38.86045,
    37.83053, 37.0899,
  77.70703, 75.72316, 70.61813, 68.313, 69.13135, 68.94763, 70.09106,
    71.94067, 74.40459, 74.99821, 74.51194, 75.21438, 75.41212, 74.42829,
    72.4318, 70.66109, 67.96465, 64.21166, 60.702, 57.35474, 54.2571,
    51.5731, 48.71611, 47.13713, 47.05245, 46.2704, 43.59927, 40.27473,
    38.85698, 37.69786,
  76.53975, 72.717, 66.76756, 63.9416, 64.16972, 64.0093, 66.41843, 70.86485,
    74.46628, 74.26525, 73.31914, 74.35139, 75.01552, 74.70737, 72.93359,
    71.47715, 69.02767, 65.84402, 63.8582, 61.08971, 57.31215, 53.88137,
    50.09642, 47.91798, 47.70945, 47.03173, 45.45776, 41.83721, 39.37049,
    38.32202,
  74.98386, 71.89525, 66.47752, 62.62946, 61.78858, 61.17622, 64.12843,
    68.95108, 72.32715, 71.66715, 72.40288, 73.4305, 74.30856, 74.04504,
    72.11334, 70.2787, 67.9321, 65.52536, 63.78198, 61.61496, 58.77413,
    55.71269, 51.96857, 49.42593, 49.16018, 47.99439, 46.5663, 43.03514,
    39.06301, 37.85672,
  72.08803, 69.56293, 64.74551, 61.006, 60.2664, 58.59194, 60.11719,
    62.64597, 64.45972, 64.64529, 66.31535, 68.2821, 70.29018, 70.47343,
    68.97198, 67.49537, 65.14454, 62.9217, 61.82086, 60.12127, 57.76802,
    55.40479, 52.74052, 51.06123, 50.64989, 49.79126, 49.04509, 46.11434,
    40.59167, 37.62504,
  66.03016, 63.91344, 60.66047, 58.56879, 59.00626, 58.01729, 56.895,
    56.27737, 55.40625, 55.47582, 55.78873, 57.67433, 59.9974, 60.68369,
    60.53476, 60.01292, 58.03346, 56.61717, 56.29262, 56.06055, 54.28513,
    51.63339, 48.56687, 47.27147, 47.61442, 47.30316, 46.76718, 46.00401,
    43.46115, 38.85583,
  50.01173, 50.78795, 51.24046, 51.73628, 53.16396, 54.80241, 52.20794,
    48.4498, 47.32088, 47.50797, 46.91043, 46.58026, 46.46207, 46.61745,
    46.53363, 46.69615, 46.26255, 45.47063, 45.02171, 44.6112, 44.69953,
    44.59407, 43.74195, 42.78524, 42.99828, 43.24503, 42.57943, 40.92244,
    40.28524, 38.98495,
  43.46943, 43.83202, 43.9369, 43.72306, 44.63643, 46.83001, 47.39467,
    43.8599, 42.03224, 43.05368, 43.52805, 43.68062, 43.11217, 42.25114,
    41.8682, 41.72765, 40.5822, 39.38462, 39.13384, 39.17017, 38.93069,
    39.46699, 40.04148, 40.22428, 40.26463, 40.53064, 40.24414, 38.99261,
    37.99031, 37.19577,
  47.50349, 47.49942, 47.37085, 47.45243, 47.33826, 47.48893, 47.75309,
    47.91429, 48.0653, 48.49377, 49.34091, 48.88852, 46.45272, 45.94106,
    45.38828, 44.27047, 43.37193, 42.72739, 42.03032, 41.84319, 41.35349,
    39.93454, 40.06504, 41.38397, 42.1075, 40.72224, 41.66944, 42.76727,
    34.48603, 31.68711,
  52.23866, 52.03833, 51.13938, 51.30456, 50.76971, 50.63665, 51.12934,
    51.61226, 51.95546, 51.94708, 52.08126, 52.29275, 52.36448, 52.05574,
    51.88501, 52.0112, 51.84544, 51.87295, 51.86483, 51.85275, 51.70202,
    51.17913, 50.85294, 51.92277, 52.15226, 46.9967, 38.2113, 40.62875,
    34.55891, 32.39147,
  54.20853, 54.05212, 53.79667, 53.48269, 53.11736, 52.8065, 52.56102,
    52.40692, 52.17887, 52.05001, 52.08844, 52.26538, 52.49432, 52.80764,
    52.9539, 52.65987, 52.61099, 52.72552, 52.84369, 52.97211, 53.33339,
    53.56653, 53.55462, 53.63871, 53.19161, 51.71109, 47.63295, 40.06142,
    34.0786, 32.79264,
  54.84985, 54.59746, 54.42459, 54.20425, 54.02623, 53.93225, 53.7386,
    53.40443, 53.0877, 52.80532, 52.75261, 53.06401, 53.22113, 53.033,
    53.49743, 53.68307, 52.99317, 52.53198, 52.92221, 53.41002, 53.9135,
    53.93256, 54.0923, 54.75504, 54.33048, 53.05645, 51.52086, 47.2419,
    37.45863, 32.61922,
  55.45428, 55.03588, 54.88743, 54.50784, 54.12727, 54.05216, 54.02711,
    53.74086, 53.47112, 53.17437, 53.15818, 53.85734, 54.38258, 54.34008,
    54.43374, 54.72258, 54.14925, 52.9683, 52.94079, 53.40247, 53.23642,
    52.64837, 53.014, 54.02356, 54.40608, 53.54347, 52.18782, 52.33553,
    52.02819, 40.573,
  55.7873, 55.7528, 55.6641, 55.35267, 54.61326, 54.57077, 55.09003, 54.7515,
    54.20721, 53.88163, 54.08974, 54.89447, 55.66774, 55.57001, 56.09621,
    56.58923, 55.88862, 54.44194, 53.06429, 53.2016, 52.77747, 47.96641,
    52.4337, 53.40533, 53.86559, 53.61885, 52.87304, 53.48406, 52.39828,
    36.04265,
  55.99483, 56.07213, 56.08416, 55.86591, 55.29193, 55.45456, 56.12622,
    56.03328, 55.41725, 54.88354, 54.56211, 53.98394, 53.39108, 53.76589,
    54.284, 54.7002, 54.61357, 53.62989, 52.69811, 52.91295, 52.66518,
    51.00421, 53.12162, 53.84199, 53.63441, 52.72548, 52.94069, 52.79197,
    51.05642, 30.78534,
  56.13554, 56.28014, 56.49806, 56.55471, 56.22616, 56.55568, 57.02556,
    56.00325, 55.08358, 55.00008, 54.72728, 54.53842, 54.514, 54.65128,
    54.80404, 55.14949, 55.3822, 55.06075, 54.21826, 53.7843, 53.50468,
    53.75856, 54.33614, 54.45165, 53.66282, 53.38709, 53.90107, 52.96009,
    45.45427, 31.39043,
  57.27437, 57.22223, 57.03786, 56.74846, 56.14723, 56.05948, 55.7971,
    56.43557, 56.8484, 56.93887, 56.95084, 56.88302, 57.15807, 58.20523,
    58.56031, 57.12664, 57.3971, 57.7957, 57.33455, 55.89001, 54.80439,
    55.19155, 55.77561, 54.99778, 53.88391, 54.58108, 53.85745, 52.02738,
    33.31879, 31.87483,
  58.75438, 59.33001, 58.40499, 58.27971, 57.45077, 55.96654, 54.49068,
    55.35077, 55.58608, 56.17611, 56.48984, 56.7064, 56.3848, 56.0408,
    55.56993, 56.61733, 57.15318, 57.21661, 57.05868, 57.1259, 57.16086,
    55.55954, 53.8772, 52.28172, 52.86392, 53.68674, 52.26721, 39.57817,
    31.29913, 30.28742,
  59.07542, 58.63324, 59.49503, 58.16703, 58.79132, 56.81625, 55.69821,
    55.37165, 55.86166, 56.51554, 54.76459, 50.58233, 48.20917, 48.33665,
    47.99012, 49.36666, 50.99017, 52.29136, 53.60408, 54.51141, 56.12934,
    54.74574, 51.92561, 51.14003, 51.63232, 51.40081, 39.15804, 31.74359,
    32.07951, 30.47146,
  64.00271, 61.51574, 63.12101, 63.63868, 61.32761, 58.92942, 56.85405,
    54.56543, 52.97618, 53.06511, 52.86259, 52.42363, 52.82024, 53.17358,
    49.49122, 49.40261, 48.4698, 48.39176, 48.63904, 51.17386, 54.49487,
    54.17892, 51.65117, 52.0505, 51.91339, 49.29177, 32.0201, 35.74008,
    32.92595, 31.39428,
  62.7257, 64.09673, 65.51274, 66.57672, 66.09158, 63.68296, 57.45305,
    54.13824, 55.73467, 54.28712, 54.60866, 54.61435, 55.36158, 55.40617,
    53.63134, 52.54646, 52.66754, 52.73979, 52.42974, 52.90152, 53.85529,
    53.18549, 49.35899, 44.94182, 43.82626, 40.24678, 33.00123, 34.48079,
    34.22429, 32.41711,
  55.51837, 55.86111, 56.18496, 55.43845, 55.2763, 55.6573, 56.51567,
    56.7869, 54.94474, 55.7467, 56.56837, 56.83146, 58.35241, 57.59637,
    55.94049, 53.86406, 52.97828, 53.3768, 53.6993, 53.37058, 52.84589,
    49.659, 43.12989, 36.7177, 33.3693, 33.07457, 31.90523, 31.5017,
    32.00242, 31.68297,
  57.63535, 57.67057, 56.74063, 55.81292, 55.1888, 55.6195, 57.33361,
    57.40892, 55.38718, 55.43979, 55.4701, 54.76062, 55.0393, 55.88958,
    55.27236, 53.6931, 53.25434, 53.59355, 54.21173, 53.57127, 44.26375,
    41.63921, 36.34953, 34.54018, 34.42068, 33.28033, 32.11677, 31.51643,
    31.02218, 30.74513,
  58.19741, 58.8226, 58.71899, 58.00828, 57.46627, 57.81558, 58.2296,
    57.34961, 55.82994, 54.53763, 54.27121, 53.62249, 53.2521, 54.09412,
    53.49756, 52.8993, 53.12513, 52.65002, 50.35914, 45.66721, 38.28648,
    38.17699, 34.89479, 33.92471, 33.97022, 33.22103, 31.97547, 31.62245,
    31.25033, 30.83304,
  57.06235, 56.76385, 56.69069, 56.83367, 56.97482, 56.80916, 57.05687,
    57.70407, 57.37482, 56.25672, 54.96768, 55.58393, 56.79499, 55.68195,
    54.09341, 53.63291, 53.21702, 51.6271, 51.0083, 46.82649, 38.57991,
    38.69424, 35.74484, 34.07102, 33.77152, 33.38863, 31.71473, 30.8122,
    30.81591, 30.70129,
  57.08779, 56.59126, 55.44901, 55.98845, 55.93509, 56.00498, 56.35535,
    57.04023, 57.48272, 57.06185, 57.64061, 58.29913, 58.25106, 58.0699,
    56.91005, 56.42628, 56.24261, 56.5136, 55.87866, 51.70617, 40.87832,
    38.66344, 36.30986, 35.01714, 33.47327, 32.66159, 31.95479, 30.58444,
    30.54962, 30.48207,
  66.84377, 62.40282, 54.47549, 50.66998, 52.46841, 53.00746, 54.76678,
    55.66098, 55.72832, 56.04406, 56.65277, 56.42014, 55.56448, 55.90075,
    55.87362, 56.81805, 59.06262, 60.98069, 60.44501, 58.13558, 50.50651,
    42.55341, 38.38461, 36.33694, 34.0806, 32.68094, 31.84399, 30.86501,
    30.53561, 30.50662,
  66.58093, 62.06858, 54.35239, 49.87327, 50.7806, 51.02793, 51.89825,
    52.99764, 54.81785, 55.64895, 55.51283, 52.97089, 53.18867, 51.8494,
    50.16414, 49.54954, 52.48343, 56.89458, 57.67631, 57.25769, 53.70984,
    47.2657, 41.4202, 38.56607, 36.1489, 33.48534, 32.08261, 31.00973,
    30.52239, 30.48687,
  67.21259, 63.53743, 55.72807, 51.34707, 51.11197, 50.67719, 50.93722,
    51.55618, 53.01332, 54.2753, 51.79842, 48.89913, 51.37402, 51.05505,
    49.26066, 48.08232, 48.3894, 49.23387, 50.28275, 49.43938, 48.75042,
    48.77026, 45.74954, 41.84967, 38.32386, 34.67542, 32.3229, 31.08149,
    30.47619, 30.49963,
  68.52897, 66.12601, 61.07072, 57.39479, 57.23802, 55.4407, 55.08666,
    54.82817, 56.2787, 55.98441, 51.53459, 49.16822, 50.22123, 49.77032,
    48.52385, 47.92241, 47.15873, 47.15259, 47.45484, 47.4571, 47.35049,
    46.30725, 46.00315, 45.21334, 41.64555, 36.1138, 33.00815, 31.84324,
    30.69021, 30.44434,
  69.86279, 68.70417, 64.06306, 61.88979, 62.34508, 61.98391, 61.38395,
    60.84634, 61.08586, 60.50126, 56.60789, 56.8219, 56.80583, 56.13959,
    54.14563, 53.04426, 51.45279, 48.66344, 47.06427, 46.22147, 45.56926,
    44.34997, 43.14079, 44.07174, 44.89808, 40.30333, 35.16077, 33.37437,
    31.8926, 30.62913,
  70.36719, 69.10845, 65.45355, 63.48166, 63.45892, 62.96689, 63.25702,
    63.98634, 65.95144, 66.00497, 65.27868, 66.31358, 67.15989, 67.17838,
    66.03558, 64.78729, 61.86915, 57.50804, 52.90539, 50.21006, 48.38885,
    46.66312, 44.55073, 43.84591, 45.08286, 45.41108, 41.13421, 35.61143,
    33.70036, 31.58735,
  70.31123, 67.88164, 63.51997, 61.2359, 60.94967, 60.73174, 62.04412,
    64.86603, 67.69128, 66.86224, 65.91179, 66.99723, 68.02871, 68.25999,
    67.23819, 66.65351, 64.99338, 61.98135, 59.234, 56.07484, 53.07342,
    50.02591, 46.44555, 44.26841, 44.55674, 45.22532, 44.25074, 39.05605,
    35.33397, 33.21248,
  70.244, 67.66036, 63.52511, 60.77676, 60.13365, 59.89317, 61.8068,
    65.09332, 66.86349, 65.62222, 65.99075, 66.9574, 68.02167, 67.74139,
    66.33365, 65.81053, 64.89159, 63.20259, 61.77058, 59.90358, 57.89214,
    55.48139, 51.33697, 48.26181, 47.82547, 46.67993, 45.80627, 40.87234,
    33.93661, 32.18599,
  67.94335, 65.3766, 61.90793, 59.68253, 59.44185, 58.77237, 60.23198,
    62.35563, 63.4235, 63.19376, 63.99654, 65.14915, 66.52477, 66.78609,
    65.8717, 65.01556, 63.45016, 62.09208, 61.18211, 59.8969, 58.58106,
    58.07163, 56.6474, 54.57493, 53.96444, 53.24083, 52.91611, 48.46386,
    37.08211, 31.11503,
  62.99111, 61.33376, 59.01328, 57.89287, 58.54128, 58.37832, 58.51536,
    58.74413, 55.93253, 56.53359, 57.3987, 59.18775, 60.90363, 61.30781,
    61.06015, 59.78344, 57.41705, 56.24804, 56.67107, 56.88126, 54.38815,
    50.78362, 47.70189, 47.00967, 48.12401, 48.50575, 48.88276, 49.785,
    44.89182, 34.20052,
  53.90439, 53.6898, 53.61625, 53.96534, 55.16523, 56.30869, 55.77419,
    51.77104, 48.90722, 49.6275, 48.94025, 48.8707, 49.30573, 49.45823,
    49.38701, 49.1544, 47.74854, 46.29903, 44.7526, 42.77069, 42.17844,
    41.60792, 39.83259, 38.50889, 39.50785, 40.35793, 39.77626, 37.73065,
    37.18472, 34.79855,
  45.67716, 46.23992, 46.07825, 45.52504, 47.58754, 52.81069, 54.6344,
    46.07654, 42.12566, 44.28256, 45.7729, 47.13514, 46.94944, 45.35104,
    43.80567, 42.52451, 39.31695, 36.02527, 35.49928, 34.99316, 33.98009,
    34.44373, 34.74274, 34.94267, 35.33677, 36.11915, 35.99887, 33.97211,
    32.00781, 30.5136,
  34.39386, 34.40742, 34.45674, 34.56916, 34.42394, 34.57346, 34.89698,
    35.3829, 36.04857, 36.96679, 39.01646, 39.03788, 35.52035, 35.88635,
    36.08277, 35.32313, 35.46733, 36.32084, 37.38019, 39.20624, 39.96129,
    38.66827, 39.4339, 42.00068, 44.12919, 44.06434, 48.97009, 51.03818,
    36.24586, 32.3756,
  38.3972, 38.6327, 37.60344, 38.30084, 37.54076, 37.1822, 37.69451,
    38.26839, 38.91639, 39.70565, 41.03476, 42.9324, 44.0233, 41.63132,
    39.76607, 40.56654, 39.53043, 40.57524, 42.28609, 43.74945, 43.49304,
    42.76429, 43.32427, 47.02694, 50.4535, 46.7196, 44.33099, 48.85702,
    37.18742, 33.68665,
  37.89339, 38.37836, 38.93062, 39.44845, 39.88209, 40.24633, 40.35722,
    40.74157, 41.2836, 41.89177, 42.62377, 44.00499, 45.3644, 47.13366,
    47.8975, 45.60597, 46.12321, 47.65701, 48.58136, 50.46498, 53.98213,
    57.46071, 58.54938, 59.19051, 58.76234, 53.8918, 51.14258, 47.18696,
    36.7774, 34.70604,
  40.71762, 41.24299, 42.58553, 43.98705, 45.31895, 46.58343, 46.47048,
    45.98133, 46.49764, 47.32818, 47.79471, 48.56878, 48.13133, 46.98665,
    50.31364, 52.52374, 49.63267, 47.11654, 49.78796, 53.1847, 57.75499,
    58.21958, 56.93736, 62.25709, 62.67414, 60.50902, 55.4984, 46.6573,
    37.83076, 33.08312,
  43.24014, 42.5182, 44.2257, 45.50027, 46.57014, 46.92244, 46.90668,
    46.88302, 48.16379, 49.28522, 49.77724, 52.06321, 53.22289, 53.66683,
    54.73801, 56.73416, 54.90759, 49.70149, 51.04597, 55.82085, 55.358,
    49.0634, 50.82132, 57.46145, 63.43508, 60.94299, 52.61317, 56.04166,
    53.67595, 38.66927,
  45.55815, 47.61588, 51.14753, 54.32291, 54.26244, 54.68312, 57.07611,
    57.45589, 56.78943, 57.58727, 59.80166, 64.34277, 66.37972, 67.72122,
    69.56432, 71.75447, 72.79141, 64.87697, 56.05011, 56.24871, 51.78674,
    46.37556, 50.04753, 55.52295, 61.81636, 60.44401, 54.7742, 62.47684,
    58.31141, 36.91995,
  47.58975, 50.02938, 52.9282, 55.70194, 56.20747, 57.36323, 60.01677,
    61.95025, 62.40812, 61.58446, 60.74256, 57.33615, 52.83595, 55.46931,
    57.97139, 59.81517, 61.84562, 57.96001, 50.47325, 51.65181, 49.52924,
    48.83645, 52.23875, 58.39913, 59.42982, 53.1061, 53.68935, 57.55706,
    50.8067, 32.64833,
  48.48257, 50.61684, 53.99091, 56.78528, 56.55221, 59.57018, 61.10371,
    54.12414, 48.764, 50.02936, 49.54879, 49.47823, 50.11332, 53.27442,
    56.17195, 59.069, 62.57264, 61.90121, 55.75292, 54.22677, 53.26698,
    55.32836, 60.86795, 64.12518, 59.81606, 57.35311, 62.38159, 61.13694,
    48.8046, 33.20568,
  56.94246, 57.67062, 58.43441, 58.88788, 58.60025, 60.11295, 57.3486,
    57.78566, 61.15213, 63.84066, 65.86319, 68.0388, 69.48017, 72.89979,
    75.52589, 74.28017, 76.35042, 78.86212, 79.45596, 71.62986, 65.31036,
    70.85591, 79.23587, 76.69525, 66.24752, 71.43645, 69.54591, 57.95312,
    37.90124, 32.76009,
  60.5871, 61.72744, 61.49867, 62.41841, 61.98355, 61.29457, 61.01493,
    62.87311, 64.48256, 67.02617, 70.14116, 72.94366, 73.58321, 72.94102,
    71.9434, 74.20907, 76.41325, 78.28413, 79.33257, 80.85656, 81.72434,
    79.43944, 74.13739, 65.49511, 64.1766, 66.32001, 59.31464, 42.03956,
    32.59202, 30.02803,
  59.81112, 58.63638, 60.00747, 60.62265, 63.36566, 65.43134, 66.38393,
    67.48925, 69.4455, 71.02227, 66.56123, 50.82093, 49.47301, 49.51613,
    50.2658, 52.04269, 55.4784, 58.20595, 61.922, 66.68419, 73.16857,
    69.97339, 52.83207, 48.31943, 51.14519, 48.84279, 39.00017, 32.97199,
    32.22161, 30.21825,
  62.78997, 59.48931, 62.27923, 63.21249, 63.54956, 64.63103, 66.38409,
    62.83047, 56.54116, 50.95694, 47.4833, 45.55334, 48.02335, 49.548,
    48.98284, 48.57668, 47.50372, 48.23574, 49.77388, 55.66231, 66.88348,
    64.87061, 48.92527, 55.58412, 55.88292, 43.97477, 33.32928, 35.08596,
    33.4362, 31.3663,
  65.68565, 66.65832, 68.37984, 68.92507, 69.20341, 67.83983, 63.45675,
    63.8243, 66.36119, 59.36563, 57.2476, 55.0259, 58.85236, 62.1655,
    60.03329, 52.50443, 53.98825, 54.86553, 59.2034, 67.07331, 64.09126,
    58.44349, 48.89243, 46.25213, 45.24943, 40.1417, 33.9446, 34.77635,
    34.81794, 32.36913,
  58.08033, 58.49044, 59.43185, 60.04612, 60.6582, 60.80577, 62.24771,
    64.26842, 63.75978, 65.26385, 67.64063, 67.95801, 70.04614, 71.49257,
    70.50529, 61.102, 58.19374, 61.56597, 65.19834, 63.36565, 55.44007,
    49.89716, 45.97168, 39.5452, 36.16592, 35.0351, 32.91164, 32.31018,
    32.63395, 31.75602,
  54.84458, 55.52468, 56.54963, 57.74906, 59.2364, 60.8316, 63.80985,
    66.2864, 66.42371, 67.92445, 67.78387, 63.79923, 67.91971, 70.13773,
    68.24901, 67.81137, 63.80224, 63.38452, 67.60153, 64.66415, 45.11338,
    44.09217, 38.97305, 37.66472, 36.8043, 34.85194, 33.16482, 31.97799,
    31.22828, 30.65976,
  55.68681, 56.7809, 58.47897, 59.82326, 61.33772, 64.00687, 67.13696,
    68.50021, 67.0211, 63.10411, 64.40037, 59.67968, 56.49289, 62.55925,
    60.11722, 59.36031, 61.02687, 57.76518, 58.20404, 53.84335, 39.73305,
    40.83567, 37.09517, 36.23752, 36.296, 35.06723, 32.81773, 32.31514,
    31.57184, 30.77694,
  54.39633, 52.84227, 54.71151, 56.81998, 59.11891, 60.70761, 63.95068,
    65.94769, 67.67849, 66.35699, 60.40305, 65.6429, 73.23759, 69.66509,
    59.90344, 57.857, 55.26438, 54.11811, 57.46828, 54.57138, 39.05238,
    40.91888, 37.87894, 36.27508, 35.76004, 35.12495, 32.52234, 31.03779,
    30.92492, 30.64304,
  51.36188, 52.36481, 52.30304, 54.70967, 57.21374, 58.60712, 60.78982,
    62.97041, 62.68718, 62.38795, 69.2944, 72.67307, 73.87, 73.74951,
    71.70254, 65.66258, 57.30618, 57.53542, 62.78336, 54.10975, 40.06817,
    39.20292, 37.27919, 36.61496, 34.34934, 33.17805, 32.49342, 30.45257,
    30.43767, 30.24338,
  57.66202, 54.57034, 49.77695, 47.68076, 49.31276, 49.73545, 50.53483,
    51.54175, 51.43457, 53.98554, 59.83894, 58.90512, 51.7453, 56.38807,
    60.21189, 64.3553, 74.29585, 79.72824, 76.71573, 68.87725, 49.98793,
    42.0712, 38.40645, 36.5752, 33.80305, 32.38442, 31.83583, 30.75731,
    30.37476, 30.23197,
  55.64967, 53.52037, 49.36184, 44.7886, 46.01099, 46.81849, 48.1839,
    49.73933, 52.37829, 59.66523, 62.02476, 53.44235, 52.76492, 51.72676,
    50.81385, 51.7323, 57.73968, 63.42091, 62.69148, 64.15874, 56.4744,
    48.14031, 41.44327, 38.61942, 36.13694, 33.06245, 31.80827, 30.79715,
    30.31866, 30.22231,
  52.90873, 51.4171, 47.63758, 44.42629, 44.56429, 44.87507, 45.27094,
    46.4363, 49.64862, 54.20444, 51.73565, 46.0968, 49.94449, 49.25229,
    47.01105, 44.57729, 44.95309, 46.27873, 49.07555, 49.76217, 50.18851,
    52.4875, 48.24342, 43.59814, 39.08165, 34.67741, 32.07775, 30.98724,
    30.3538, 30.23542,
  52.84538, 48.55676, 45.78622, 44.13466, 44.34713, 43.01909, 43.97058,
    44.95028, 49.39399, 51.58905, 45.01484, 40.45683, 43.57534, 44.44605,
    44.11247, 44.50608, 44.64133, 45.36847, 46.81889, 47.26517, 47.49786,
    48.58347, 50.09196, 49.35884, 43.37711, 36.16187, 32.44315, 31.60763,
    30.60319, 30.2079,
  53.34755, 52.57842, 48.35259, 46.30658, 49.54084, 50.77762, 49.78119,
    47.58838, 49.19221, 47.90739, 41.57113, 42.06305, 43.50611, 44.9943,
    44.60701, 45.76796, 46.02891, 43.73698, 42.89771, 42.70483, 42.21442,
    42.26656, 42.11345, 44.26697, 46.70239, 41.12607, 34.9347, 33.58785,
    32.08306, 30.35714,
  57.30136, 56.86887, 55.32501, 53.40871, 54.59914, 53.75102, 55.7649,
    56.77116, 59.22516, 53.73272, 45.72779, 47.79737, 49.72904, 51.58812,
    51.35346, 51.70215, 52.13807, 49.91365, 46.11172, 44.56875, 43.13703,
    42.04795, 41.42018, 41.2755, 43.57276, 45.81242, 41.51801, 35.6502,
    33.81379, 31.29075,
  61.61288, 59.10196, 52.48932, 50.67325, 52.35862, 52.34949, 52.67702,
    55.72015, 60.79019, 56.15568, 48.73808, 51.5256, 51.73876, 52.95765,
    53.52333, 55.29728, 55.38329, 54.86907, 51.9539, 48.24144, 46.38974,
    45.11275, 43.74461, 42.72761, 44.10605, 47.56826, 47.37334, 41.61261,
    37.48242, 33.97938,
  63.29861, 61.79284, 60.29288, 54.66673, 53.14506, 52.75654, 56.81785,
    61.19887, 59.34705, 53.98138, 53.48258, 54.9198, 54.56847, 53.97915,
    52.79456, 54.79227, 56.77143, 57.52941, 56.2766, 52.92218, 50.97404,
    49.86406, 46.45171, 43.24092, 44.07217, 46.0032, 48.22387, 44.14352,
    35.99441, 33.22147,
  64.07627, 61.56228, 60.09719, 55.7456, 54.5408, 52.18725, 56.5414,
    58.50227, 54.82653, 53.30441, 55.44527, 55.13651, 54.62062, 54.79688,
    55.62769, 57.69783, 59.94374, 62.07954, 62.07868, 60.04044, 59.44426,
    61.84941, 62.43978, 58.81122, 56.16361, 56.07588, 58.78414, 54.49291,
    39.24331, 30.9618,
  62.77607, 60.34901, 60.23483, 60.32508, 61.93685, 62.75714, 61.44541,
    57.15283, 50.54361, 52.54281, 53.37636, 53.94046, 54.339, 54.97572,
    57.41241, 58.76163, 58.98236, 60.46495, 62.12628, 63.27331, 60.19227,
    56.51988, 53.589, 52.92849, 53.54422, 54.83683, 56.38781, 59.38378,
    52.65129, 35.39874,
  55.28696, 55.80697, 57.28999, 59.0621, 60.70831, 62.22699, 62.27912,
    55.31912, 50.81549, 51.79866, 51.38588, 52.70595, 54.08124, 54.55496,
    56.00914, 56.30259, 54.49101, 52.67484, 49.2285, 44.91365, 43.72612,
    42.18623, 39.53204, 38.05546, 39.77428, 41.82953, 42.56292, 41.18338,
    40.94113, 36.80069,
  54.04055, 57.14793, 57.68334, 53.71226, 59.48604, 64.63821, 66.12701,
    57.62508, 50.94914, 54.5183, 57.2211, 61.15633, 61.6176, 57.57592,
    54.38179, 52.48394, 47.03614, 40.90854, 39.61694, 37.67887, 35.38785,
    35.32609, 35.15519, 35.20516, 35.86644, 37.24723, 37.6615, 35.39481,
    32.49696, 30.25479,
  31.16283, 31.43532, 31.73144, 32.05892, 32.23901, 32.50886, 32.85605,
    33.27906, 33.78214, 34.43328, 35.96539, 36.00791, 34.03309, 34.47475,
    34.70466, 34.2765, 34.48441, 35.05745, 35.74503, 37.08924, 37.89766,
    37.62033, 38.39353, 39.7352, 40.55262, 40.32601, 43.59186, 43.64516,
    34.29673, 31.35228,
  35.60402, 36.14105, 35.97537, 36.89068, 36.98827, 37.22543, 37.86525,
    38.5667, 39.33929, 40.15528, 41.16333, 42.48512, 43.21449, 41.81168,
    41.0847, 41.55038, 40.99112, 41.66952, 42.79181, 43.71084, 43.66039,
    43.32711, 43.94451, 46.8363, 50.46027, 48.50325, 45.34554, 45.90538,
    35.45013, 32.3824,
  37.81065, 38.57027, 39.30808, 40.19909, 41.02863, 41.91549, 42.7563,
    43.7868, 44.90272, 45.92057, 46.97042, 48.36198, 49.59822, 51.20741,
    52.0779, 51.04996, 51.54731, 52.42696, 52.61972, 53.54223, 55.30374,
    56.89606, 57.24485, 57.90632, 59.0512, 56.37277, 51.05178, 44.80058,
    35.72421, 33.36106,
  43.09389, 44.62397, 46.32671, 48.11149, 49.87658, 51.79504, 52.90852,
    53.77615, 55.22264, 56.62188, 57.38943, 58.29486, 58.65891, 58.74711,
    61.12932, 62.61208, 60.66435, 58.38649, 58.98274, 59.93367, 62.39124,
    61.49985, 58.44979, 63.0618, 64.43691, 58.91617, 53.8609, 43.33083,
    35.49191, 31.91938,
  48.48692, 49.46482, 51.27909, 53.04314, 54.54894, 55.68265, 56.74285,
    58.07819, 60.19574, 61.62138, 61.6516, 62.00516, 62.45504, 63.45095,
    64.10398, 64.29546, 62.29836, 58.57717, 58.39696, 62.95789, 64.05757,
    56.52373, 56.20282, 58.97194, 61.95757, 59.03072, 51.77808, 51.4532,
    46.79287, 35.22981,
  53.87189, 56.54261, 59.35436, 62.27549, 63.14708, 63.65707, 65.52889,
    67.13207, 68.39599, 70.41298, 72.4566, 75.1855, 75.64199, 75.16035,
    75.10735, 76.04435, 77.0046, 73.57912, 63.63407, 62.87591, 58.53698,
    53.98198, 54.76303, 56.17001, 58.89443, 57.07586, 53.81915, 61.37952,
    54.53501, 33.84779,
  63.91199, 67.61095, 70.54884, 73.42477, 74.50346, 74.75745, 75.44554,
    75.50605, 74.96086, 74.64114, 74.47082, 70.69624, 65.79398, 64.90128,
    67.48997, 72.02946, 70.88052, 63.68205, 57.88325, 56.99268, 54.50139,
    52.84372, 53.53543, 55.98123, 56.00869, 52.68941, 54.43612, 59.54562,
    49.61962, 31.30855,
  68.67909, 71.29723, 72.98795, 74.19206, 73.03562, 73.80721, 73.4201,
    65.94962, 61.17605, 60.38639, 59.06335, 57.75311, 56.92513, 57.805,
    59.64242, 61.17942, 61.55907, 59.75622, 55.07608, 53.94718, 52.64899,
    52.58756, 54.71102, 56.13711, 53.52256, 52.65792, 58.73964, 56.86186,
    41.87687, 31.74136,
  71.27737, 72.27312, 72.89896, 72.13225, 70.51781, 70.47901, 66.95034,
    65.84887, 68.03194, 69.60379, 70.67165, 71.82404, 73.2915, 78.71797,
    79.34049, 73.92819, 72.71658, 73.81921, 71.60049, 65.97064, 62.50373,
    65.51189, 70.02877, 67.34425, 59.46951, 60.03853, 59.32255, 49.98551,
    35.70264, 31.4647,
  78.55407, 80.12242, 81.02607, 82.14555, 81.60062, 80.10916, 79.66918,
    80.62645, 81.15488, 81.89425, 82.38349, 83.10324, 82.88033, 81.60293,
    80.24378, 80.60101, 80.62071, 78.95234, 72.22266, 68.3377, 67.70707,
    64.81853, 61.92971, 56.47528, 59.30044, 67.39513, 55.38977, 36.80451,
    31.6757, 29.96918,
  80.8581, 82.06322, 84.0905, 84.99535, 86.8212, 85.95172, 84.73662,
    84.22986, 83.92342, 84.45455, 84.13872, 79.25394, 78.48623, 77.07278,
    74.94375, 72.86377, 70.93826, 67.36803, 62.8609, 59.68595, 60.29665,
    55.48306, 47.35714, 43.15684, 44.09642, 43.10145, 36.2816, 31.38372,
    30.84278, 29.90181,
  82.85051, 79.83689, 82.93505, 84.93638, 85.1025, 84.08645, 83.39098,
    80.84397, 78.05808, 77.67644, 75.02399, 69.60578, 70.17778, 69.97845,
    66.00638, 62.75534, 58.91338, 56.17775, 53.38086, 52.15686, 52.95191,
    48.2945, 40.7952, 45.62893, 47.67229, 36.31421, 31.17961, 31.84152,
    31.29122, 30.36886,
  87.52453, 87.95898, 89.71606, 90.73769, 90.07635, 87.30399, 80.88344,
    77.49487, 78.14183, 76.08516, 76.64456, 76.01109, 76.18581, 76.37193,
    70.94673, 61.95021, 59.73886, 56.60697, 54.10419, 55.00853, 52.82418,
    45.35579, 41.41794, 42.08386, 42.1945, 34.50305, 31.82248, 32.06968,
    32.06489, 30.8909,
  83.82602, 84.48783, 84.5709, 82.91357, 81.54253, 80.64745, 80.4529,
    80.96387, 78.76439, 78.8158, 79.61828, 77.97757, 79.09222, 79.59324,
    77.68327, 76.06796, 69.93825, 69.27608, 67.61425, 62.42834, 51.75569,
    45.51952, 44.88987, 37.41239, 33.78423, 32.90764, 31.61026, 31.05996,
    31.2285, 30.67085,
  76.94042, 77.04491, 76.79748, 76.3923, 76.34391, 77.66863, 81.66841,
    83.0331, 80.45706, 80.57433, 80.38519, 79.91696, 79.79119, 78.86614,
    77.7067, 76.02912, 73.73071, 67.34988, 65.95169, 60.81308, 46.51708,
    42.85728, 36.68629, 34.26289, 32.99623, 32.48699, 31.52095, 30.87716,
    30.53952, 30.19868,
  77.07011, 77.9466, 78.62782, 78.9038, 79.15657, 80.48465, 81.82172,
    81.98355, 81.59555, 80.63734, 80.022, 78.44889, 77.53577, 77.77762,
    76.357, 70.811, 65.8873, 57.71767, 53.92095, 49.3752, 38.56464, 37.49364,
    34.88328, 34.0068, 33.29179, 32.41488, 31.53397, 31.05337, 30.66856,
    30.20069,
  77.34141, 77.78768, 78.23797, 78.69831, 79.5013, 79.65319, 80.33576,
    81.15907, 80.73003, 79.87815, 78.43869, 78.54704, 79.44577, 77.65189,
    69.33096, 63.67178, 57.91836, 52.20669, 52.31731, 49.53128, 37.15528,
    37.19702, 35.31345, 34.11891, 33.037, 32.41878, 31.40018, 30.55097,
    30.41009, 30.16799,
  74.13363, 76.00549, 76.94911, 77.54076, 77.84666, 78.44576, 78.79221,
    79.33208, 79.77812, 78.78347, 78.73018, 79.02846, 78.23009, 76.16449,
    73.44176, 63.14591, 52.68984, 48.04863, 50.22853, 46.63472, 37.60571,
    36.74216, 34.94851, 33.76799, 32.07665, 31.64484, 31.19652, 30.22369,
    30.10929, 29.96186,
  71.61002, 71.03335, 69.44846, 69.28022, 70.54884, 71.24541, 72.79411,
    74.12763, 73.23482, 72.7378, 74.3934, 71.46701, 65.50711, 66.89838,
    66.96046, 64.5845, 63.55639, 63.13156, 63.49202, 57.15228, 45.03591,
    38.23495, 34.91071, 33.58809, 31.67518, 31.071, 30.78261, 30.26672,
    30.04165, 29.92727,
  66.43591, 65.67535, 64.59003, 63.65417, 64.53219, 65.59778, 67.14075,
    68.33792, 69.24023, 71.77645, 71.04299, 64.58244, 63.67146, 64.11749,
    63.45763, 61.64264, 61.42181, 61.14198, 59.66659, 56.70142, 49.29846,
    41.33686, 35.83909, 34.14857, 32.39056, 31.26029, 30.72606, 30.28759,
    30.02285, 29.93574,
  61.43256, 61.08554, 60.27046, 59.89919, 60.57468, 61.74719, 63.18348,
    64.44964, 65.77965, 67.04729, 63.36578, 58.33176, 59.22604, 58.48119,
    56.22917, 53.20383, 51.50594, 50.2612, 50.03837, 48.52293, 46.19557,
    44.15734, 39.72182, 36.04543, 33.50858, 31.86072, 30.75517, 30.32094,
    30.04033, 29.94368,
  60.53518, 57.49392, 56.81351, 56.7302, 57.46934, 57.62446, 58.50515,
    58.70295, 60.1458, 59.37114, 53.88948, 50.9128, 51.24082, 50.04335,
    48.34065, 46.8779, 45.33535, 44.25331, 43.64454, 42.72955, 43.29358,
    43.83602, 42.4176, 41.29867, 37.03005, 32.83507, 30.98808, 30.6075,
    30.10717, 29.94507,
  58.15066, 56.17776, 54.5352, 54.3485, 56.0848, 56.77614, 55.77354,
    53.72636, 53.50209, 51.06667, 46.5578, 46.35831, 46.57857, 46.28126,
    45.31648, 45.01197, 44.13533, 41.93181, 40.67727, 40.00776, 40.72135,
    41.28555, 39.38591, 39.63078, 39.2198, 35.13065, 31.80748, 31.45952,
    30.66125, 30.00398,
  62.02138, 60.3284, 59.81178, 59.84702, 60.072, 59.53582, 59.71575,
    58.67165, 57.47467, 52.29696, 48.2116, 49.73315, 50.37381, 50.36451,
    49.27417, 47.91933, 46.70278, 44.36766, 41.45972, 40.49377, 40.80761,
    40.43641, 38.74536, 37.76232, 38.07877, 37.96388, 34.80248, 32.12291,
    31.28934, 30.32728,
  65.80066, 67.70094, 63.72964, 62.965, 63.68813, 63.03387, 61.03157,
    59.99706, 60.57154, 56.71872, 52.03621, 53.69741, 53.99771, 53.05636,
    51.32491, 49.84632, 47.60639, 45.72306, 42.93477, 40.44779, 40.37125,
    39.93716, 38.38887, 37.00929, 36.07337, 37.09182, 37.04354, 34.37113,
    32.9449, 31.3918,
  73.84572, 77.79768, 74.80134, 71.13277, 68.9708, 67.05804, 66.80994,
    65.65311, 61.57493, 57.46193, 55.69235, 56.32352, 56.00805, 53.28078,
    50.27052, 48.77226, 47.27477, 45.78444, 43.63369, 41.11743, 41.02073,
    40.81655, 38.5154, 36.63208, 36.1932, 36.44775, 37.48117, 35.86137,
    32.63896, 31.15192,
  77.19386, 79.19251, 74.04212, 71.08083, 69.47971, 67.11034, 66.70379,
    63.91743, 58.39647, 55.8525, 55.9842, 56.00019, 54.89204, 52.4483,
    50.46408, 49.02548, 47.77457, 47.03915, 45.57223, 43.99708, 45.24709,
    47.14466, 46.16887, 42.65284, 40.27704, 39.72257, 40.79992, 39.5552,
    33.40713, 30.1972,
  76.02881, 76.67348, 74.20172, 73.81496, 73.44076, 70.48537, 67.57147,
    62.51981, 56.85294, 56.74303, 56.71131, 57.04723, 56.60802, 55.24572,
    54.60309, 53.49035, 51.95178, 51.38631, 50.9278, 50.69379, 51.15619,
    49.82247, 46.26436, 43.69239, 42.0153, 41.41837, 40.83303, 42.27738,
    39.17474, 31.93337,
  70.77987, 71.52528, 75.16466, 77.98224, 77.62425, 76.16732, 70.59165,
    62.55209, 59.33329, 59.70303, 58.87716, 58.69283, 58.88785, 59.49769,
    60.05495, 59.23185, 57.56404, 55.52802, 51.69613, 47.76783, 46.20363,
    44.1769, 41.61567, 39.78435, 39.30199, 39.00992, 38.08057, 36.44455,
    35.79821, 32.96044,
  70.02553, 72.05803, 73.38426, 73.72525, 74.03207, 76.02368, 74.31231,
    66.01297, 62.13605, 63.93394, 64.75189, 65.12699, 64.24097, 62.80811,
    60.70451, 57.1062, 51.80573, 46.34961, 43.57039, 40.97835, 38.93304,
    37.88398, 36.88004, 36.07116, 35.54574, 35.4804, 34.89212, 33.23033,
    31.57161, 30.20617,
  31.9023, 31.98001, 32.06186, 32.14374, 32.15584, 32.19921, 32.2682,
    32.37489, 32.5619, 32.79185, 33.71217, 33.84535, 32.50166, 32.68547,
    32.82531, 32.48853, 32.4472, 32.64268, 32.86958, 33.5726, 34.03594,
    33.59484, 33.7688, 34.6895, 35.50583, 35.46966, 38.15785, 39.52998,
    34.3927, 32.71472,
  32.85739, 33.01567, 32.73841, 33.10261, 32.96988, 32.88506, 33.06533,
    33.2535, 33.49105, 33.76111, 34.15108, 34.77976, 35.16505, 34.33084,
    33.87293, 34.18338, 33.84321, 34.23614, 35.03518, 35.79145, 35.97197,
    35.95069, 36.62921, 38.19961, 42.73088, 43.74965, 39.0215, 41.11694,
    35.06421, 33.30049,
  32.81182, 32.90837, 32.97614, 33.10817, 33.21984, 33.35428, 33.52187,
    33.7678, 34.03329, 34.27235, 34.58215, 35.18538, 35.6777, 36.47224,
    37.05918, 36.57608, 37.08248, 38.02192, 38.57768, 39.52913, 41.24831,
    43.29705, 44.46841, 44.13068, 47.95269, 50.05882, 42.05561, 40.27683,
    35.02398, 33.91711,
  33.85907, 34.1711, 34.67939, 35.22634, 35.81195, 36.5979, 36.88614,
    36.86203, 37.26608, 37.88876, 38.31342, 38.966, 39.25101, 39.26944,
    41.10659, 42.9119, 42.52906, 41.68606, 42.73596, 43.97757, 46.70203,
    47.7167, 45.79968, 50.50915, 52.54302, 46.04576, 44.8428, 39.296,
    34.97585, 33.03508,
  37.03883, 37.2049, 37.93464, 38.67125, 39.18975, 39.49704, 39.77773,
    40.00328, 40.84483, 41.58836, 41.69477, 42.145, 42.72523, 43.74342,
    44.88951, 46.02099, 45.61316, 44.3726, 44.8131, 49.93501, 51.78736,
    43.84923, 43.85899, 45.32424, 46.9446, 45.44234, 41.4645, 41.32068,
    40.64252, 35.08794,
  40.25855, 41.13489, 42.38993, 43.84035, 43.78441, 43.49082, 44.25728,
    44.78901, 45.0777, 45.98759, 47.23343, 50.04428, 53.04262, 53.06944,
    52.73473, 61.51874, 70.86584, 57.00667, 47.54882, 48.19437, 45.56047,
    41.93303, 42.6144, 43.71467, 45.83002, 44.37872, 47.01535, 61.54652,
    53.4981, 34.04649,
  44.68975, 46.25491, 47.96059, 49.8158, 50.7077, 51.485, 53.30075, 55.49634,
    55.7722, 55.43115, 55.3616, 53.72484, 51.2495, 51.03037, 55.58287,
    61.81362, 57.14607, 49.00798, 45.32094, 44.67774, 43.05417, 42.03847,
    42.7207, 44.95129, 45.62506, 42.12183, 50.953, 66.72227, 51.45499,
    32.41215,
  50.46072, 52.50251, 54.38295, 56.15131, 56.25626, 57.83832, 59.13953,
    55.0033, 51.60078, 50.64015, 49.11162, 47.17848, 45.58464, 45.51959,
    46.43627, 47.35257, 47.18038, 46.07464, 43.28585, 42.52169, 41.59729,
    41.34017, 42.79337, 44.54941, 43.49831, 41.49477, 52.55306, 57.70395,
    39.33665, 33.07076,
  56.33771, 57.13329, 57.79926, 57.27379, 55.88751, 55.53134, 52.23251,
    49.66777, 49.44406, 48.87438, 47.86311, 47.02981, 46.74605, 50.52409,
    52.98575, 47.91148, 47.41842, 48.80507, 48.23238, 44.96124, 42.60194,
    44.78097, 49.04121, 49.10587, 44.49387, 45.10067, 48.52494, 45.27875,
    35.55588, 32.95955,
  61.5514, 63.58719, 63.12601, 62.93107, 60.21756, 54.66925, 49.14161,
    50.2533, 50.82135, 52.52103, 54.72971, 58.46412, 58.65309, 55.47208,
    52.00224, 53.1624, 54.21082, 53.71939, 51.30304, 49.79738, 50.24482,
    49.83647, 49.13536, 45.52357, 52.83086, 66.01342, 52.6326, 36.32073,
    33.27719, 31.94954,
  78.91154, 78.75951, 78.79268, 75.57007, 74.24202, 68.8905, 64.56477,
    66.53692, 67.24709, 75.57949, 80.6319, 56.62107, 52.11348, 51.42511,
    51.452, 52.05172, 52.78006, 52.07495, 50.49352, 49.59171, 51.28106,
    49.14071, 43.91533, 40.4753, 42.3828, 43.80442, 37.6418, 32.89283,
    32.44656, 31.83623,
  84.62353, 80.58965, 83.45175, 84.40247, 83.94466, 82.59312, 81.56274,
    74.567, 64.01759, 63.90807, 60.95789, 52.42729, 54.27641, 54.50481,
    51.04718, 51.099, 49.45849, 48.25637, 46.75647, 46.04033, 47.17924,
    44.74935, 38.83395, 42.79212, 45.10006, 35.51575, 32.49968, 32.91333,
    32.68044, 32.10714,
  91.10452, 91.39768, 94.30395, 94.39257, 92.81814, 88.49792, 80.7327,
    71.7021, 71.27106, 64.41116, 63.88725, 58.31673, 60.22372, 60.82279,
    53.77495, 49.77595, 48.24972, 46.55113, 44.93475, 45.87607, 45.64417,
    41.33781, 37.86004, 41.44628, 43.17691, 34.44669, 32.93192, 33.12413,
    33.23857, 32.48736,
  90.01748, 92.76633, 91.53619, 88.33717, 85.18419, 82.88914, 81.7465,
    81.32148, 78.51497, 77.46675, 78.46082, 77.04823, 77.94902, 78.17383,
    75.06741, 58.69099, 49.08349, 50.15309, 50.16708, 48.94266, 43.71389,
    42.42846, 45.17673, 38.28073, 34.93246, 33.81324, 32.96103, 32.61027,
    32.77732, 32.37666,
  81.96161, 81.38495, 79.83656, 78.08459, 76.64614, 78.25185, 83.83719,
    83.57386, 79.84711, 78.93315, 77.84348, 72.92017, 64.83424, 68.76247,
    70.17117, 54.79171, 53.35477, 50.98853, 51.53508, 52.28684, 48.12547,
    41.7921, 36.5631, 34.59179, 33.6838, 33.70565, 32.95927, 32.46006,
    32.27909, 32.04901,
  77.52713, 77.20756, 77.13934, 76.59173, 76.21967, 77.02837, 77.95896,
    77.58804, 73.73786, 69.26399, 65.86253, 60.33986, 56.6259, 57.87951,
    54.93786, 52.04889, 50.93416, 47.03879, 45.76826, 44.28075, 38.19827,
    36.2949, 34.25137, 33.87827, 33.88736, 33.56594, 32.95452, 32.5435,
    32.2721, 31.99992,
  72.02161, 70.49224, 69.59391, 69.0303, 68.90982, 67.91844, 67.11093,
    66.16903, 63.85659, 61.53216, 57.03814, 56.80186, 59.29668, 54.78899,
    50.90741, 48.69843, 46.26893, 43.19622, 43.76235, 42.63223, 35.41504,
    35.59897, 34.67637, 33.93966, 33.62352, 33.52443, 32.9012, 32.28862,
    32.15919, 32.00034,
  64.82351, 64.44395, 62.88232, 61.97087, 60.5775, 59.96384, 59.19473,
    58.41732, 57.89938, 55.31154, 55.4336, 56.91578, 54.68183, 52.79276,
    52.57969, 48.27304, 42.82809, 39.99582, 42.06618, 40.93656, 35.56137,
    35.51087, 34.75884, 34.08047, 33.19715, 33.06571, 32.76557, 32.09542,
    31.99129, 31.89858,
  62.57591, 61.0082, 57.77873, 55.4981, 54.62632, 53.56791, 53.04586,
    52.81386, 51.65663, 50.61402, 51.67153, 49.90642, 45.21314, 45.51495,
    45.80552, 44.94009, 45.15838, 45.92947, 48.10522, 46.76957, 40.75656,
    36.87704, 34.70671, 34.15439, 33.00955, 32.66687, 32.49492, 32.10606,
    31.95452, 31.87019,
  58.38116, 56.36388, 53.3249, 50.73309, 49.92332, 49.154, 48.56095,
    47.92149, 47.34336, 48.70697, 48.38191, 43.81604, 42.82818, 43.48919,
    43.86335, 43.68899, 44.8457, 46.30808, 47.28128, 47.18655, 43.61238,
    38.64397, 35.04885, 34.43087, 33.44587, 32.73674, 32.40854, 32.13017,
    31.94492, 31.86895,
  53.97747, 52.19338, 49.46874, 47.25618, 46.30399, 45.71577, 45.18192,
    44.79173, 45.19709, 46.65786, 44.84899, 41.81207, 43.31635, 44.1517,
    43.93984, 42.96035, 42.54768, 42.11497, 42.17313, 41.44878, 40.03108,
    39.00242, 37.07303, 35.36881, 34.01754, 33.0947, 32.44969, 32.14189,
    31.96368, 31.87739,
  52.6559, 49.78808, 47.5054, 45.85215, 45.08578, 44.13451, 43.99342,
    43.77674, 45.25839, 46.00704, 43.02435, 41.27466, 42.30515, 42.36262,
    41.71062, 40.85217, 39.68447, 38.71542, 38.19353, 37.3893, 38.49951,
    39.51048, 37.80855, 38.08314, 36.00661, 33.68395, 32.5571, 32.29723,
    32.00089, 31.88849,
  51.33768, 49.50198, 47.06706, 45.66645, 46.04079, 46.19822, 45.4931,
    44.16358, 44.44518, 43.31801, 40.11904, 39.6268, 39.8884, 39.90483,
    39.24874, 38.99175, 38.44901, 37.13293, 36.49473, 36.07457, 37.24397,
    38.0108, 35.9292, 36.91827, 37.12967, 34.86654, 32.92291, 32.79757,
    32.35626, 31.93964,
  52.01995, 50.64943, 49.49293, 48.7859, 48.32998, 47.4145, 47.06682,
    46.33602, 45.95208, 42.39688, 38.7539, 39.17117, 39.66872, 40.19128,
    39.99223, 39.54351, 39.28697, 38.27983, 36.7187, 36.10917, 36.26139,
    36.15328, 35.4417, 35.33329, 35.98045, 36.22419, 34.61452, 33.18938,
    32.71252, 32.11407,
  52.16566, 52.43984, 49.53535, 48.17316, 47.95934, 47.03938, 45.46089,
    44.64017, 45.25473, 42.30318, 38.35351, 39.25223, 40.16591, 40.65646,
    40.5705, 40.40768, 39.65255, 39.11288, 37.80756, 36.32695, 36.27568,
    36.32193, 35.91118, 35.15561, 34.62961, 35.68231, 35.84175, 34.30256,
    33.64186, 32.74152,
  52.94611, 54.39351, 52.54073, 49.69797, 47.72556, 46.22948, 46.29982,
    46.40721, 44.41721, 41.30001, 39.61067, 40.43417, 41.43044, 41.11443,
    40.21112, 39.98267, 39.54388, 39.13645, 38.26735, 36.75951, 36.6662,
    36.78291, 35.64895, 34.70832, 34.65041, 35.09064, 36.11321, 35.30653,
    33.50922, 32.56627,
  53.48676, 54.07877, 50.7782, 48.28946, 46.97936, 45.49784, 46.07126,
    45.55185, 42.3987, 40.26652, 40.26794, 40.82402, 41.14931, 40.61918,
    40.13791, 39.69413, 39.12136, 38.9016, 38.11847, 36.83007, 37.27485,
    38.61097, 38.74452, 37.44818, 36.73637, 36.82964, 37.99711, 37.66373,
    33.97537, 31.96151,
  52.49759, 51.65842, 49.37661, 48.63556, 48.35781, 47.08258, 46.50346,
    44.3103, 40.61044, 40.10421, 39.91463, 40.23463, 40.49414, 40.37077,
    40.61164, 40.21911, 39.4101, 39.37458, 39.53057, 39.62561, 40.3086,
    40.34273, 39.137, 38.15627, 37.64581, 37.70576, 37.72433, 39.10265,
    37.34948, 33.01136,
  49.88873, 48.55622, 48.87637, 49.44326, 49.33285, 49.44727, 47.08318,
    42.26086, 39.59218, 39.30571, 38.43534, 38.41484, 39.01676, 40.13944,
    41.60135, 42.29239, 42.37112, 42.48295, 41.34329, 39.68877, 39.30701,
    38.55811, 37.3926, 36.64631, 36.64512, 36.80574, 36.53871, 35.8708,
    35.73534, 33.73343,
  49.49905, 49.24988, 48.80823, 47.88399, 47.42014, 49.0169, 48.88567,
    43.72747, 40.54629, 41.1949, 41.83136, 42.85862, 43.58904, 44.26083,
    44.69566, 44.2949, 42.56135, 40.30625, 39.09435, 37.76393, 36.74974,
    36.25872, 35.797, 35.4135, 35.17977, 35.30985, 34.99335, 34.01669,
    33.1347, 32.16445,
  29.16066, 29.20716, 29.25703, 29.29981, 29.2784, 29.27961, 29.30096,
    29.33982, 29.43878, 29.57193, 30.27543, 30.41671, 29.46916, 29.60529,
    29.72588, 29.4288, 29.3315, 29.40414, 29.48281, 29.97424, 30.26682,
    29.80967, 29.78217, 30.36883, 30.83786, 30.71003, 33.03008, 34.46048,
    30.94107, 29.80929,
  29.66391, 29.77178, 29.56481, 29.8183, 29.67916, 29.5427, 29.63168,
    29.72691, 29.86941, 30.05758, 30.36263, 30.84293, 31.17802, 30.54414,
    30.08506, 30.19846, 29.78571, 29.89956, 30.37374, 30.87646, 30.90272,
    30.59878, 30.88597, 31.8648, 35.79173, 37.17459, 33.67896, 35.91254,
    31.5011, 30.22924,
  29.71806, 29.73778, 29.71966, 29.76379, 29.75953, 29.7998, 29.84385,
    29.95751, 30.08076, 30.17406, 30.32366, 30.7009, 30.96502, 31.36473,
    31.54638, 30.86016, 30.89356, 31.38577, 31.62018, 32.14475, 33.28227,
    34.73932, 35.76783, 35.44074, 40.02253, 43.22375, 35.868, 35.37328,
    31.40327, 30.68085,
  30.05473, 30.12341, 30.34474, 30.59183, 30.87122, 31.31207, 31.42696,
    31.27484, 31.41044, 31.70529, 31.86336, 32.23202, 32.19006, 31.85295,
    32.92308, 34.03179, 33.58843, 32.82893, 33.54238, 34.48945, 36.93866,
    38.257, 36.87606, 41.49876, 44.13058, 38.85756, 38.30802, 34.61837,
    31.45103, 30.06221,
  31.36165, 31.22175, 31.60465, 32.02357, 32.31997, 32.4651, 32.54456,
    32.53167, 32.97612, 33.31282, 33.15028, 33.25149, 33.43258, 33.92481,
    34.73858, 35.57517, 35.17561, 34.76439, 35.4477, 40.44812, 42.73249,
    36.235, 36.20086, 37.71082, 39.28672, 38.13986, 35.49992, 35.2405,
    35.30257, 31.60739,
  32.65422, 33.02186, 33.79235, 34.73526, 34.53332, 34.04676, 34.32205,
    34.42343, 34.35438, 34.74191, 35.34293, 37.36655, 39.72839, 40.00186,
    39.49578, 47.76747, 57.68444, 46.54462, 38.67092, 40.08566, 38.32669,
    34.97258, 35.36809, 36.02048, 37.87015, 36.96857, 39.36606, 52.70884,
    47.49195, 30.85465,
  34.43573, 35.11134, 36.0231, 37.04582, 37.34549, 37.65336, 38.9384,
    40.7647, 41.48214, 41.88573, 42.61704, 42.20088, 40.92769, 40.87996,
    46.16591, 54.08314, 49.83608, 40.96628, 37.85546, 37.35048, 35.8709,
    34.93569, 35.36823, 37.17926, 38.14768, 35.2268, 44.32454, 61.13502,
    47.34967, 29.5154,
  36.95632, 38.16571, 39.6042, 41.22412, 41.80715, 43.83296, 46.07434,
    44.18734, 42.58146, 42.61834, 41.99564, 40.65375, 39.26865, 38.95855,
    39.97445, 40.94514, 39.68361, 38.24635, 36.26088, 35.73902, 35.01673,
    34.68087, 35.86486, 37.46216, 36.86905, 34.71524, 46.38326, 53.23474,
    35.51965, 30.42223,
  42.32571, 43.56363, 44.96985, 45.61776, 45.74127, 46.68011, 45.06759,
    43.49196, 43.30476, 42.79046, 41.67487, 40.37918, 39.49791, 42.07037,
    43.59252, 39.23773, 38.71082, 39.88093, 39.55204, 37.11849, 35.13242,
    36.56971, 40.04522, 40.36615, 36.7372, 37.23476, 41.68333, 40.63515,
    32.82314, 30.38795,
  48.60497, 51.24817, 51.90862, 52.41993, 51.08191, 47.10408, 42.5524,
    42.62411, 42.34728, 42.61839, 43.69641, 46.79567, 47.23581, 44.94091,
    41.98087, 41.98061, 42.48098, 42.16129, 40.7341, 40.15348, 40.48462,
    40.85515, 41.13483, 38.82013, 44.66144, 55.53309, 46.37615, 33.49911,
    30.88525, 29.36405,
  70.9642, 73.90285, 66.34411, 56.79553, 55.31805, 52.19597, 48.1473,
    50.26013, 51.6939, 60.27926, 67.76035, 47.48805, 42.12654, 40.85074,
    40.0758, 40.22206, 41.03761, 41.5083, 40.22581, 39.92763, 42.49233,
    41.8596, 37.9878, 35.2768, 38.30888, 41.13339, 35.38739, 30.33009,
    29.77427, 29.20423,
  79.53227, 74.55636, 77.11783, 78.31673, 77.55126, 65.96396, 66.106,
    60.20937, 50.74918, 53.64967, 53.12975, 41.21175, 42.45045, 42.87785,
    39.63308, 40.49591, 39.36064, 38.99541, 38.17482, 38.35973, 40.88252,
    39.39294, 34.32585, 37.68559, 39.79463, 32.43266, 29.64756, 30.09021,
    29.96093, 29.41371,
  82.03358, 81.99027, 86.95467, 88.09747, 88.48228, 85.63267, 75.12733,
    52.4385, 52.80376, 48.54796, 47.02657, 42.15047, 45.44745, 46.92615,
    41.19498, 40.40913, 39.78761, 38.64667, 37.56698, 39.36683, 40.47527,
    36.73302, 33.43861, 37.79551, 39.55358, 31.40698, 29.94536, 30.21902,
    30.4645, 29.76964,
  84.39507, 90.10918, 89.29165, 87.06667, 84.22075, 80.61582, 76.93477,
    76.50473, 69.44374, 65.14904, 73.38549, 69.94292, 71.7729, 70.31602,
    60.56068, 47.66205, 40.06345, 41.65997, 42.91417, 43.36889, 39.2591,
    37.75734, 39.80211, 34.88527, 32.26313, 30.74402, 30.03127, 29.77043,
    30.08455, 29.69879,
  76.73105, 76.84247, 71.33767, 66.67879, 61.78106, 71.27188, 79.37885,
    79.94253, 77.31161, 76.71246, 76.20521, 61.27533, 50.35291, 55.82241,
    60.2154, 44.4694, 44.26207, 43.59863, 46.5955, 47.91583, 42.52141,
    37.90044, 33.74829, 31.43093, 30.48256, 30.7699, 30.11806, 29.67719,
    29.58506, 29.39016,
  60.71022, 58.42995, 57.13732, 55.86632, 56.30359, 60.70727, 65.54655,
    63.50459, 60.63121, 57.29839, 53.09941, 47.22736, 44.3105, 46.89199,
    46.0804, 43.54766, 44.26658, 41.83929, 42.13615, 41.62653, 35.3403,
    32.75892, 30.75159, 30.63452, 30.87429, 30.68458, 30.16824, 29.77835,
    29.58681, 29.33748,
  55.8381, 54.19591, 53.51186, 53.50683, 54.11284, 53.97868, 53.45214,
    52.96412, 51.35725, 48.96851, 45.11681, 45.70695, 49.24847, 46.15799,
    43.2104, 42.32962, 40.8304, 38.47313, 39.94029, 39.13186, 31.65721,
    31.7757, 31.28303, 30.79072, 30.6386, 30.6548, 30.13377, 29.5459,
    29.48541, 29.34367,
  52.19794, 52.15402, 51.43647, 51.20675, 50.43261, 49.87812, 49.3272,
    48.81221, 47.65441, 45.4465, 45.82267, 48.16396, 46.8408, 45.40583,
    46.26254, 43.03373, 37.94911, 35.21761, 38.09551, 37.46019, 31.89732,
    32.10927, 31.66659, 31.10357, 30.297, 30.29716, 30.01756, 29.37651,
    29.30627, 29.24369,
  52.51578, 51.73466, 49.40605, 47.6811, 46.83519, 45.94849, 45.6278,
    45.52541, 44.59177, 43.86387, 45.65214, 44.63943, 39.69633, 39.57793,
    39.83602, 38.69076, 38.51268, 38.94184, 41.69151, 41.06833, 35.66168,
    33.18449, 31.88231, 31.27979, 30.18025, 29.93756, 29.78683, 29.38825,
    29.27563, 29.21777,
  50.92628, 49.45885, 46.98155, 44.9229, 44.30572, 43.90554, 43.61452,
    43.25484, 42.82507, 44.34839, 44.34819, 39.25902, 36.57704, 36.25905,
    35.91247, 35.26869, 36.61665, 38.65679, 40.80476, 41.84029, 38.99405,
    35.05949, 32.24102, 31.50261, 30.55766, 29.97527, 29.72089, 29.4377,
    29.28193, 29.21322,
  48.21014, 47.19567, 45.31635, 43.447, 42.82338, 42.42777, 41.94011,
    41.3401, 41.32779, 42.60088, 40.095, 35.52326, 35.67236, 35.91291,
    35.58378, 34.81108, 35.00906, 35.47417, 36.74022, 37.11617, 36.29856,
    35.62056, 34.00327, 32.19129, 31.00412, 30.28637, 29.71957, 29.43422,
    29.29245, 29.22334,
  47.3377, 46.0492, 44.03791, 42.5926, 41.81335, 40.67975, 40.10057,
    39.35033, 40.31459, 40.71277, 37.11478, 34.58194, 35.23352, 35.32936,
    34.95952, 34.55233, 34.01884, 33.66018, 33.65484, 33.14212, 34.23403,
    35.25903, 34.70195, 35.06321, 33.14017, 30.93285, 29.8121, 29.56621,
    29.31426, 29.2245,
  45.52937, 44.99783, 42.47307, 40.97946, 41.12808, 41.01279, 40.13782,
    38.9413, 39.67893, 38.81731, 35.39434, 34.56096, 34.73424, 34.67887,
    34.10166, 34.09101, 33.81863, 32.7185, 32.14027, 31.85869, 33.24495,
    33.86287, 32.57314, 34.07058, 34.44762, 32.04226, 30.09076, 30.05571,
    29.63653, 29.27475,
  45.10246, 43.68002, 42.50623, 41.83715, 41.57729, 41.09652, 41.29877,
    41.52271, 42.38913, 39.36966, 35.25214, 35.17379, 35.26228, 35.44177,
    35.05574, 34.71115, 34.6503, 33.71176, 32.33048, 31.96244, 32.42318,
    32.45028, 31.88644, 32.13346, 33.22864, 33.51004, 31.75576, 30.41708,
    30.01667, 29.4466,
  44.29842, 44.64935, 42.06902, 41.10072, 41.4888, 41.37739, 40.81713,
    41.12911, 42.83706, 39.8762, 35.23521, 35.32772, 35.60414, 35.59824,
    35.31359, 35.25269, 34.81053, 34.54681, 33.34085, 31.9496, 32.21194,
    32.55886, 32.40491, 31.71574, 31.1902, 32.42661, 32.6394, 31.25737,
    30.87127, 30.00502,
  44.92477, 46.69584, 45.48072, 43.44568, 42.03085, 41.06264, 42.07038,
    43.28269, 41.88616, 38.40963, 35.79574, 35.85024, 36.3541, 35.62065,
    34.65024, 34.61904, 34.49186, 34.52587, 33.76932, 32.28179, 32.65728,
    33.11152, 32.04239, 31.14622, 30.93115, 31.48138, 32.79869, 32.16753,
    30.76956, 29.85597,
  46.39639, 47.6721, 44.71544, 42.67441, 41.60364, 40.52684, 41.91193,
    42.42878, 39.41301, 36.70069, 35.991, 36.00889, 35.89521, 35.04278,
    34.52251, 34.2732, 34.04594, 34.2747, 33.63644, 32.20113, 32.90903,
    34.60916, 34.86589, 33.45617, 32.61832, 32.8574, 34.54688, 34.51963,
    31.10747, 29.28241,
  45.93277, 45.63934, 43.52335, 42.83501, 42.9556, 42.16236, 42.32163,
    40.79702, 37.089, 36.20017, 35.6584, 35.59821, 35.43268, 34.83577,
    34.93024, 34.63756, 33.93808, 34.01434, 34.1418, 34.07623, 35.47187,
    36.30628, 35.26826, 33.93189, 33.20984, 33.45651, 33.84828, 35.85316,
    34.34595, 30.22433,
  43.29948, 42.05, 42.37826, 43.51862, 44.25416, 45.14769, 43.48464,
    39.24328, 36.60435, 36.12999, 34.78948, 33.91457, 33.59431, 33.9693,
    35.06457, 35.70549, 35.93895, 36.44496, 35.52909, 34.08809, 34.22412,
    33.83522, 32.73011, 32.04816, 32.1652, 32.62887, 32.75133, 32.64132,
    33.05566, 30.94717,
  42.34741, 42.19035, 42.11658, 41.81535, 41.95595, 44.34797, 44.92271,
    40.00344, 36.68777, 36.78107, 36.61386, 36.59973, 36.40433, 36.89055,
    37.69197, 37.66925, 36.5124, 34.95227, 33.95025, 32.68831, 31.94607,
    31.63815, 31.39896, 31.22879, 31.26167, 31.68517, 31.67777, 31.01976,
    30.4233, 29.53295,
  22.43003, 22.46362, 22.5019, 22.53378, 22.51888, 22.50551, 22.50373,
    22.53289, 22.59198, 22.69338, 23.53358, 23.68184, 22.69496, 22.84762,
    22.95997, 22.63785, 22.56243, 22.61769, 22.65248, 23.1953, 23.50214,
    22.97466, 22.89097, 23.39199, 23.71036, 23.44229, 26.00471, 27.79601,
    24.43238, 23.18059,
  22.85246, 22.91291, 22.68215, 22.93966, 22.76624, 22.60374, 22.66829,
    22.73139, 22.84132, 23.02104, 23.40577, 23.99007, 24.37351, 23.68203,
    23.1973, 23.27508, 22.81884, 22.87729, 23.36206, 23.89226, 23.81576,
    23.27683, 23.30775, 24.1904, 27.9279, 28.78682, 26.68728, 29.8161,
    25.22808, 23.73236,
  22.7888, 22.80752, 22.76172, 22.79054, 22.75166, 22.73957, 22.76164,
    22.8433, 22.96097, 23.05404, 23.16949, 23.59304, 23.93285, 24.3579,
    24.4292, 23.59088, 23.52892, 23.9309, 24.01244, 24.28083, 25.15428,
    26.59468, 27.54892, 27.15697, 31.66835, 34.47634, 29.02276, 29.31903,
    25.10574, 24.32451,
  22.85561, 22.87793, 23.05022, 23.21111, 23.45866, 23.89692, 23.97376,
    23.80532, 23.88693, 24.15114, 24.31486, 24.68268, 24.49776, 24.09286,
    25.07648, 26.07111, 25.4744, 24.44276, 24.76608, 25.35105, 27.92115,
    29.40226, 28.29419, 32.76088, 34.91869, 31.29337, 31.7873, 28.57648,
    25.1642, 23.58728,
  23.59044, 23.33012, 23.61559, 23.95107, 24.22131, 24.41399, 24.45667,
    24.38948, 24.86001, 25.2377, 25.09425, 25.05633, 24.9064, 25.20165,
    25.98894, 26.67498, 26.02203, 25.28566, 25.92703, 30.7152, 32.70638,
    27.50068, 27.32922, 29.25915, 31.12238, 30.43387, 28.57015, 28.81932,
    29.28544, 25.18658,
  24.12651, 24.29645, 25.03612, 26.02994, 25.90577, 25.3941, 25.56629,
    25.42974, 25.0687, 25.1549, 25.37439, 27.28122, 29.63413, 29.73617,
    29.29282, 36.49635, 44.31641, 35.55137, 29.39778, 31.41076, 29.69544,
    26.14204, 26.58185, 27.42117, 29.85722, 29.28263, 31.03419, 43.24813,
    39.66213, 24.60912,
  25.34519, 25.76805, 26.5328, 27.4526, 27.55365, 27.38238, 28.22354,
    29.75752, 30.1135, 30.22323, 30.97648, 30.74622, 29.69231, 29.9279,
    35.73, 43.51987, 40.13727, 31.98559, 29.03312, 28.78064, 27.19339,
    26.05667, 26.53819, 28.83554, 30.25909, 27.57608, 36.59514, 52.77948,
    40.59267, 23.16586,
  27.00093, 27.58186, 28.62227, 29.77232, 29.89564, 32.00912, 34.50653,
    32.52187, 30.89301, 31.06735, 30.72264, 29.48982, 28.30394, 28.46665,
    30.58726, 32.29776, 30.92258, 29.39585, 27.46823, 27.00773, 26.28941,
    25.86745, 27.21317, 29.57205, 29.18701, 27.31434, 39.80942, 46.66692,
    29.91859, 23.46984,
  30.70875, 31.28491, 32.57999, 33.07943, 33.47694, 35.29997, 34.2901,
    32.6798, 32.61879, 32.33974, 31.08711, 29.49779, 28.52997, 31.78348,
    33.89523, 29.81919, 29.51829, 30.99871, 30.88244, 28.4506, 26.16855,
    27.57048, 31.81828, 32.78313, 29.06274, 29.59971, 36.15601, 34.9845,
    25.60174, 23.48753,
  35.91251, 38.28214, 40.12647, 41.80589, 41.18684, 37.37388, 32.99449,
    32.88403, 32.24941, 31.63518, 32.17882, 35.40919, 36.54698, 34.89714,
    32.35499, 32.25072, 32.99453, 33.35046, 31.72248, 29.87943, 29.95023,
    30.55687, 31.55415, 29.91711, 35.06725, 45.78994, 38.81252, 26.73079,
    23.97825, 22.68274,
  51.95932, 55.49378, 50.65245, 44.09726, 42.46614, 40.90272, 36.89507,
    38.82848, 40.5136, 47.88705, 52.68435, 37.04727, 31.86707, 30.6192,
    29.63099, 30.30553, 31.32961, 31.09205, 29.86072, 29.60011, 32.08247,
    31.62269, 28.79293, 26.78399, 30.74041, 34.81184, 29.00241, 23.43535,
    23.01021, 22.50556,
  67.87675, 55.35751, 57.11819, 58.33457, 57.09151, 49.40719, 51.34846,
    48.1456, 41.06867, 44.72256, 44.06124, 30.62794, 30.90142, 31.50496,
    29.3239, 29.66238, 28.87552, 28.50516, 28.13684, 28.90052, 31.64086,
    30.48534, 26.34665, 29.38951, 31.36418, 25.43179, 22.86948, 23.30885,
    23.20967, 22.6925,
  77.7766, 73.97273, 87.21329, 89.77414, 91.66212, 83.18352, 63.20401,
    43.67325, 42.41393, 39.25008, 36.04348, 29.26253, 33.09903, 35.43342,
    30.74306, 29.67121, 29.50505, 28.77913, 28.06507, 30.29079, 31.79881,
    28.61117, 25.75229, 30.34978, 31.91632, 24.55453, 23.13121, 23.47451,
    23.75355, 23.02791,
  83.63082, 90.97022, 91.97503, 91.39844, 81.4999, 71.37579, 68.32483,
    62.24569, 53.16892, 47.62997, 54.16024, 52.25824, 54.44405, 53.33684,
    46.33551, 36.12176, 29.81109, 31.71803, 33.08838, 34.11764, 30.98014,
    29.59158, 31.42774, 28.06998, 25.59739, 23.81931, 23.23245, 23.06547,
    23.46377, 22.9864,
  63.0105, 67.78758, 63.33319, 58.82963, 52.26071, 57.70251, 77.77559,
    75.80962, 66.54559, 66.11134, 63.27784, 50.0237, 39.81412, 44.87125,
    47.44555, 33.96842, 33.99836, 33.81982, 36.56966, 37.52946, 33.76561,
    30.34306, 27.26256, 24.64447, 23.49994, 23.88157, 23.30902, 22.93593,
    22.93538, 22.70309,
  50.26917, 48.57719, 46.78211, 44.57848, 44.08772, 48.66049, 54.63132,
    53.1323, 50.49001, 48.2948, 44.42452, 37.0072, 32.31291, 35.47353,
    35.35464, 33.50658, 34.9478, 33.18018, 33.98853, 33.82533, 28.66114,
    25.88098, 23.74529, 23.60646, 23.94199, 23.78375, 23.36553, 23.04087,
    22.8809, 22.62152,
  45.52362, 43.07579, 41.54034, 41.08494, 41.99432, 42.86094, 43.23766,
    43.19806, 41.84899, 39.37089, 34.64486, 33.3341, 36.32195, 34.70176,
    33.13189, 33.19728, 32.62517, 30.88873, 32.60077, 31.65161, 24.60621,
    24.51897, 24.19757, 23.82204, 23.76602, 23.77313, 23.30396, 22.82021,
    22.78298, 22.61452,
  40.52697, 39.88498, 39.40792, 39.94499, 40.17654, 40.61003, 40.51649,
    39.98857, 38.88442, 35.40289, 34.08516, 36.17544, 36.13877, 35.4534,
    37.01918, 34.70386, 30.46109, 27.99051, 30.97682, 30.11652, 24.58849,
    24.85816, 24.58137, 24.12307, 23.43691, 23.46992, 23.18191, 22.66521,
    22.61825, 22.52859,
  40.72549, 40.87017, 39.53077, 38.78376, 38.64482, 38.13999, 37.70263,
    37.10539, 35.48808, 33.59278, 34.90378, 34.76595, 30.95208, 31.39599,
    32.29763, 31.19372, 30.54461, 30.66353, 33.48915, 32.73815, 27.79659,
    25.82015, 24.79594, 24.32996, 23.33881, 23.14938, 23.03146, 22.66543,
    22.56449, 22.49903,
  41.36995, 41.07618, 39.23761, 37.52619, 37.10586, 36.59332, 36.11836,
    35.46355, 34.33774, 35.0432, 35.30527, 31.09021, 28.40153, 28.44679,
    28.15454, 27.28589, 28.44473, 30.41089, 32.81325, 33.91013, 31.21598,
    27.63028, 25.1685, 24.47268, 23.68396, 23.1933, 22.9784, 22.71157,
    22.57403, 22.50368,
  40.70669, 40.21802, 38.21098, 36.58965, 36.08773, 35.8789, 35.55645,
    34.86823, 34.46824, 35.36156, 32.66925, 27.76043, 27.53745, 27.75132,
    27.25215, 26.35909, 26.63881, 27.42713, 29.11776, 29.96367, 29.30258,
    28.44747, 26.84061, 25.08871, 24.05288, 23.46832, 22.9929, 22.71429,
    22.595, 22.50939,
  40.82448, 39.2655, 37.56159, 36.42503, 36.05598, 35.44952, 35.15364,
    34.29822, 34.49385, 33.91301, 29.3975, 26.24454, 26.70679, 26.81357,
    26.55161, 26.27488, 26.00075, 26.00166, 26.3327, 26.0841, 27.1123,
    27.94855, 27.69996, 27.91997, 26.15245, 24.05776, 23.08205, 22.81967,
    22.62229, 22.52846,
  39.98516, 39.005, 37.10568, 35.97541, 36.40734, 36.58595, 35.73413,
    34.08157, 33.83006, 31.66173, 27.12521, 25.82668, 26.10678, 26.24906,
    25.9453, 26.22178, 26.1959, 25.33759, 24.83151, 24.68359, 26.08665,
    26.57071, 25.84636, 27.49115, 27.60536, 25.00361, 23.31334, 23.2784,
    22.91017, 22.55564,
  39.50024, 38.58268, 37.57043, 37.11871, 37.10492, 36.71472, 36.598,
    36.03721, 35.79752, 31.56646, 26.66252, 26.47192, 26.81961, 27.22493,
    27.06059, 26.99201, 27.09879, 26.19096, 24.99617, 24.92367, 25.49079,
    25.43733, 25.0162, 25.46613, 26.59659, 26.58316, 24.80552, 23.59231,
    23.242, 22.69711,
  39.05855, 39.6129, 37.2925, 36.42553, 36.63608, 36.24744, 35.56995,
    35.4577, 36.29025, 32.13982, 26.93196, 26.99313, 27.55181, 27.74861,
    27.64278, 27.64591, 27.28288, 27.01862, 25.91972, 24.8478, 25.23141,
    25.49981, 25.31852, 24.65504, 24.35059, 25.61206, 25.62642, 24.29127,
    24.02642, 23.12978,
  38.93808, 40.70019, 39.56318, 37.82539, 36.32325, 35.37953, 36.30658,
    37.32255, 35.57388, 31.05814, 27.68882, 27.69515, 28.43088, 27.95636,
    27.14346, 27.17721, 26.99795, 27.04162, 26.31698, 25.01883, 25.5255,
    25.88749, 24.83759, 24.00201, 23.82763, 24.47989, 25.77868, 25.02592,
    23.9705, 23.03844,
  39.96285, 41.55944, 38.75467, 36.77497, 35.7317, 34.97009, 36.54454,
    37.06325, 33.36285, 29.47685, 27.99696, 27.93614, 28.06412, 27.43413,
    27.01027, 26.81764, 26.62978, 26.83467, 26.17146, 24.90164, 25.61476,
    27.00803, 27.02607, 25.84366, 25.29095, 25.56711, 27.42293, 27.19699,
    24.1119, 22.53726,
  39.27972, 39.50555, 37.39033, 36.62656, 37.11285, 36.79905, 37.35423,
    35.57255, 30.96047, 28.7804, 27.58706, 27.47978, 27.47655, 27.19559,
    27.48661, 27.19028, 26.45969, 26.46867, 26.42955, 26.28114, 27.70417,
    28.32388, 27.43094, 26.28706, 25.84653, 26.0996, 26.75841, 28.81263,
    27.00334, 23.26128,
  36.57205, 35.7909, 36.25553, 37.51862, 38.83091, 40.14964, 38.61842,
    34.13539, 30.4647, 28.77094, 26.77902, 25.83242, 25.71276, 26.29701,
    27.44232, 27.84307, 27.84143, 28.3151, 27.37655, 26.17135, 26.46198,
    26.12262, 25.12784, 24.5848, 24.79799, 25.33997, 25.54326, 25.74092,
    26.20383, 23.90384,
  35.52354, 35.71307, 35.87581, 35.91537, 36.46953, 39.17672, 39.62647,
    34.35036, 30.18994, 29.05044, 28.10611, 27.81356, 27.82341, 28.58787,
    29.41171, 29.34294, 28.32162, 27.02091, 26.04397, 24.87974, 24.2872,
    24.07665, 23.91864, 23.88367, 24.01604, 24.55003, 24.62957, 24.0382,
    23.63823, 22.819,
  16.19686, 16.23071, 16.25326, 16.27566, 16.28165, 16.26768, 16.26412,
    16.2747, 16.33774, 16.3889, 17.10432, 17.21214, 16.4013, 16.52182,
    16.6085, 16.34717, 16.2906, 16.3177, 16.32604, 16.77088, 17.01534,
    16.6024, 16.50673, 16.90153, 17.13229, 16.84669, 19.07638, 20.51718,
    17.90555, 16.83117,
  16.49307, 16.52463, 16.37123, 16.58166, 16.45279, 16.31479, 16.34827,
    16.39633, 16.4776, 16.61954, 16.96123, 17.4307, 17.71104, 17.13027,
    16.79534, 16.83437, 16.44253, 16.46454, 16.84615, 17.25342, 17.17237,
    16.67239, 16.64524, 17.29086, 20.6092, 21.1385, 20.06808, 23.09516,
    18.89351, 17.44345,
  16.4428, 16.44741, 16.41037, 16.45119, 16.41519, 16.38083, 16.38288,
    16.44621, 16.53723, 16.59799, 16.69227, 17.04715, 17.31463, 17.64618,
    17.69075, 17.0231, 16.93351, 17.21483, 17.22193, 17.33912, 17.93207,
    19.08417, 19.98207, 19.53154, 23.93473, 26.66746, 22.442, 22.82486,
    18.85868, 17.98148,
  16.43947, 16.43236, 16.58081, 16.71822, 16.94215, 17.34488, 17.36166,
    17.12014, 17.15567, 17.39443, 17.50586, 17.75885, 17.57295, 17.27966,
    18.07191, 18.89742, 18.30921, 17.36159, 17.49059, 17.77651, 20.02989,
    21.41831, 20.56951, 24.63976, 26.48652, 24.23751, 25.36307, 22.28018,
    18.80628, 17.30307,
  16.86227, 16.62126, 16.8435, 17.14399, 17.41958, 17.56989, 17.5455,
    17.41515, 17.83565, 18.17044, 18.02304, 17.92023, 17.73616, 17.94035,
    18.60205, 19.03785, 18.24164, 17.61211, 18.04286, 22.42814, 24.19426,
    19.89117, 19.78125, 21.71838, 23.38222, 23.16907, 22.26644, 22.38775,
    22.72688, 18.74797,
  16.89552, 16.9733, 17.61344, 18.53166, 18.48132, 17.99677, 18.07913,
    17.90415, 17.59231, 17.66681, 17.69261, 19.26597, 21.18085, 21.34277,
    20.69096, 26.84934, 33.21231, 25.8351, 20.99024, 23.215, 21.89467,
    18.7231, 19.20573, 19.87319, 22.15485, 21.72042, 23.8535, 35.25323,
    31.85128, 18.20482,
  17.22622, 17.53933, 18.24555, 19.10234, 19.19334, 18.85514, 19.44885,
    20.77106, 21.05162, 21.07932, 21.77323, 21.65399, 20.87908, 20.99496,
    25.67844, 32.75365, 30.76197, 23.40868, 21.05917, 20.95071, 19.58567,
    18.63992, 19.07295, 21.35184, 22.87625, 20.02752, 28.8258, 44.06054,
    32.56155, 16.88528,
  17.85655, 18.19857, 19.05689, 19.98921, 19.91205, 21.73998, 23.86672,
    22.11032, 20.82763, 21.05972, 21.10953, 20.3087, 19.47768, 19.72502,
    21.90112, 23.78111, 22.59533, 21.06697, 19.72176, 19.42821, 18.88876,
    18.59877, 19.88528, 22.32249, 22.06842, 20.20729, 32.83229, 39.18979,
    23.29156, 17.11327,
  20.1128, 20.3574, 21.41671, 21.70632, 22.12486, 23.87846, 23.07671,
    21.55319, 21.58679, 21.6029, 20.91962, 20.04361, 19.58279, 22.77972,
    24.6804, 21.32984, 21.03904, 22.53149, 22.74423, 20.67761, 18.73668,
    20.02004, 24.06372, 24.99981, 21.66141, 22.14288, 29.06153, 28.08092,
    19.19308, 17.17413,
  23.55503, 25.26315, 26.88847, 28.08653, 28.17902, 25.37718, 21.69327,
    21.52668, 21.12822, 20.52111, 21.41875, 24.79569, 26.22908, 25.76324,
    24.41966, 24.04731, 24.62868, 25.196, 23.9127, 22.27872, 22.09659,
    22.8157, 24.13936, 22.82555, 27.31024, 36.74117, 30.92912, 20.23708,
    17.69162, 16.46321,
  35.95691, 39.97815, 36.36027, 31.07206, 29.96996, 28.40595, 24.71857,
    26.27437, 27.54062, 34.30085, 38.3984, 26.61036, 23.2017, 22.56452,
    21.89214, 22.61939, 23.73165, 23.56315, 22.29984, 22.01187, 24.15069,
    24.07496, 21.59767, 19.79329, 23.91894, 28.44459, 22.93579, 17.19496,
    16.74234, 16.28528,
  50.86312, 41.21188, 42.00346, 42.59263, 40.92798, 34.87814, 37.32602,
    35.05836, 29.17649, 33.62805, 33.56896, 21.48842, 22.2996, 23.10449,
    21.54037, 21.92282, 21.21846, 20.97667, 20.59474, 21.15851, 23.80545,
    22.97964, 19.37963, 22.15129, 24.09986, 19.12869, 16.67209, 17.01654,
    16.94555, 16.45704,
  58.76697, 54.71808, 70.73421, 75.27341, 74.73621, 65.90286, 50.40668,
    32.6817, 30.93412, 29.32525, 26.37682, 19.63816, 23.9838, 26.69802,
    22.70268, 21.82236, 21.68616, 20.98753, 20.45159, 22.59524, 24.23741,
    21.51707, 18.91673, 23.60785, 25.20531, 18.29904, 16.82494, 17.17975,
    17.46455, 16.76096,
  65.07981, 86.16717, 88.09285, 82.63007, 70.99954, 61.18758, 54.36032,
    47.87323, 40.53566, 35.25313, 40.84589, 39.4296, 43.16518, 43.40213,
    36.78868, 27.69161, 22.09883, 23.47444, 24.74893, 25.97501, 23.66521,
    22.61383, 24.39587, 21.84933, 19.39642, 17.41767, 16.93335, 16.81121,
    17.2392, 16.75947,
  48.56576, 55.98261, 53.46048, 50.245, 43.67479, 46.5632, 63.03461,
    61.43142, 52.09072, 51.94071, 50.70618, 39.63586, 31.60969, 37.04102,
    38.92724, 26.38601, 25.57323, 25.52776, 28.21034, 29.47762, 26.20497,
    23.72907, 21.31768, 18.54738, 17.08004, 17.46214, 17.00513, 16.68591,
    16.73107, 16.49149,
  37.57587, 37.17126, 36.33047, 34.61135, 33.57161, 37.64537, 43.90681,
    42.12357, 39.05879, 38.0889, 35.4605, 28.11261, 23.63069, 27.71935,
    27.9482, 25.29641, 26.85609, 25.30207, 26.30882, 26.4407, 22.18478,
    19.7924, 17.60187, 17.43774, 17.63465, 17.40899, 17.05607, 16.79811,
    16.67383, 16.40788,
  35.11806, 33.57279, 31.87594, 30.93582, 31.41076, 32.40977, 32.86209,
    32.46781, 31.4878, 29.54563, 25.27084, 24.33205, 27.39311, 26.10546,
    24.92654, 25.26827, 25.17531, 23.55907, 24.76357, 23.92295, 18.31902,
    18.15022, 17.96225, 17.6823, 17.51462, 17.44747, 17.01846, 16.59592,
    16.58088, 16.40379,
  31.389, 30.29801, 29.28076, 29.55103, 29.88672, 30.61077, 30.80933,
    30.34066, 29.27694, 25.90453, 24.60881, 27.12946, 27.675, 27.25303,
    28.67999, 26.86575, 23.39865, 21.32213, 23.76268, 22.79244, 18.16872,
    18.43598, 18.26312, 17.89635, 17.2031, 17.18664, 16.90798, 16.42562,
    16.41137, 16.32235,
  30.84755, 30.53455, 29.15314, 28.61945, 28.77806, 28.68671, 28.47881,
    27.79002, 25.99821, 24.05127, 25.98557, 26.73478, 23.47677, 24.28153,
    25.21421, 24.06382, 23.35011, 23.44884, 25.75843, 24.71812, 20.7311,
    19.24857, 18.40594, 18.00634, 17.07373, 16.87996, 16.76139, 16.43425,
    16.36035, 16.29175,
  31.13616, 30.86997, 29.20449, 27.77173, 27.69002, 27.36757, 26.90112,
    26.12178, 24.97361, 26.13541, 27.26331, 23.83196, 21.49503, 21.67744,
    21.39035, 20.56503, 21.51152, 23.33375, 25.15303, 25.74858, 23.88493,
    20.98337, 18.65223, 18.05728, 17.33774, 16.908, 16.72336, 16.47501,
    16.36239, 16.29431,
  30.61286, 30.39499, 28.62526, 27.16852, 26.82682, 26.67652, 26.3779,
    25.87934, 25.81047, 27.39156, 25.63718, 21.119, 20.96401, 21.0043,
    20.33965, 19.51882, 19.76029, 20.58377, 21.89569, 22.6241, 22.56633,
    21.92605, 20.15462, 18.52979, 17.68117, 17.15634, 16.73534, 16.46726,
    16.37659, 16.29958,
  30.97161, 29.79811, 28.13115, 27.08566, 26.83198, 26.46789, 26.51389,
    26.1972, 26.84471, 26.84766, 22.897, 19.73048, 20.06536, 20.02678,
    19.64674, 19.36141, 19.15197, 19.21908, 19.65377, 19.57257, 20.60379,
    21.12238, 20.43217, 20.65954, 19.4101, 17.63852, 16.80913, 16.54814,
    16.39029, 16.30514,
  30.53269, 29.60896, 27.79304, 26.88767, 27.50042, 28.03665, 27.90088,
    26.82281, 26.87097, 25.09883, 20.77871, 19.21238, 19.3096, 19.33837,
    19.05155, 19.3246, 19.35597, 18.7174, 18.38351, 18.27391, 19.5893,
    19.75877, 18.7647, 20.39062, 20.67889, 18.38952, 16.97991, 16.95545,
    16.63661, 16.33005,
  30.05761, 29.353, 28.52507, 28.39678, 28.85769, 29.0621, 29.30662,
    28.78984, 28.4502, 24.69028, 20.11283, 19.65065, 19.90516, 20.26241,
    20.0853, 20.10668, 20.2233, 19.4074, 18.41767, 18.40778, 18.8984,
    18.71742, 18.18438, 18.64222, 19.7298, 19.74745, 18.31427, 17.30531,
    16.98354, 16.45672,
  30.14314, 30.91509, 29.00248, 28.52029, 29.05321, 28.92148, 28.43788,
    28.15732, 28.77149, 25.03893, 20.28793, 20.11059, 20.50627, 20.79436,
    20.78052, 20.76254, 20.34098, 19.95879, 19.11788, 18.39689, 18.57854,
    18.62745, 18.44707, 17.9504, 17.8726, 19.10395, 19.14639, 17.92448,
    17.74487, 16.8538,
  30.77673, 32.94741, 31.64351, 29.92498, 28.82654, 27.9466, 28.54466,
    29.30504, 28.03331, 24.12904, 20.97243, 20.74605, 21.19967, 20.91088,
    20.34854, 20.30062, 19.91065, 19.85227, 19.48515, 18.59178, 18.84872,
    19.0224, 18.18861, 17.55581, 17.46482, 18.10797, 19.40714, 18.65442,
    17.73439, 16.8027,
  31.91591, 34.03235, 31.48331, 29.23422, 28.07937, 27.16404, 28.60979,
    29.34216, 26.31385, 22.79923, 21.36712, 21.10142, 21.05578, 20.51639,
    20.13642, 19.92707, 19.60633, 19.67358, 19.38813, 18.54565, 18.90241,
    19.8703, 19.79184, 19.02662, 18.81889, 19.01955, 20.83658, 20.60459,
    17.8113, 16.34939,
  31.74766, 32.29601, 29.80893, 28.59806, 28.85166, 28.50498, 29.25452,
    28.1074, 24.32952, 22.24857, 21.11034, 20.72476, 20.48337, 20.30119,
    20.59333, 20.28253, 19.52524, 19.36247, 19.57796, 19.72443, 20.45813,
    20.67998, 20.14236, 19.48191, 19.44101, 19.54979, 20.21168, 22.10052,
    20.33278, 16.95515,
  29.15774, 28.11083, 28.18243, 29.29159, 30.47279, 31.47767, 30.41329,
    26.81134, 23.70966, 22.19273, 20.33175, 19.26847, 19.05959, 19.48422,
    20.3, 20.5287, 20.44551, 20.77437, 20.31561, 19.68487, 19.79935,
    19.43981, 18.63157, 18.19567, 18.45158, 18.92374, 19.06721, 19.31532,
    19.78669, 17.52335,
  27.60538, 27.5202, 27.77905, 28.09606, 28.63959, 30.93126, 31.29743,
    26.82075, 23.28985, 22.14536, 21.10178, 20.7087, 20.77914, 21.16489,
    21.56543, 21.70611, 21.00005, 19.96758, 19.2747, 18.49314, 17.99282,
    17.84612, 17.66159, 17.58864, 17.70304, 18.21824, 18.28548, 17.68828,
    17.36747, 16.59356,
  9.868218, 9.895164, 9.924418, 9.938376, 9.939834, 9.931024, 9.918859,
    9.929762, 9.972531, 9.99791, 10.65653, 10.69627, 10.00563, 10.16769,
    10.24987, 10.00165, 9.945618, 9.967414, 9.9681, 10.38557, 10.61655,
    10.27501, 10.18723, 10.50372, 10.61306, 10.29194, 12.50966, 13.91328,
    11.62868, 10.47219,
  10.15234, 10.15078, 10.02479, 10.22047, 10.09611, 9.971257, 9.988365,
    10.02381, 10.08904, 10.19964, 10.55593, 10.96421, 11.15875, 10.67073,
    10.44782, 10.43308, 10.05372, 10.06932, 10.42096, 10.84789, 10.81065,
    10.29101, 10.20438, 10.68571, 13.88426, 14.30304, 13.62809, 16.47026,
    12.61683, 11.08938,
  10.10813, 10.09985, 10.06251, 10.11147, 10.0491, 9.986327, 9.979595,
    10.0392, 10.13076, 10.18429, 10.24439, 10.5694, 10.83084, 11.12176,
    11.13161, 10.50812, 10.42328, 10.66966, 10.68472, 10.79181, 11.22986,
    12.11776, 12.89723, 12.40351, 16.79965, 19.3345, 15.67954, 16.14667,
    12.44821, 11.54298,
  10.05372, 10.03456, 10.18, 10.299, 10.49509, 10.85703, 10.84896, 10.60921,
    10.64632, 10.88475, 10.93033, 11.10738, 10.8883, 10.68828, 11.38174,
    12.07864, 11.53819, 10.69111, 10.68904, 10.77421, 12.86248, 14.06944,
    13.35576, 17.22235, 18.92039, 17.31498, 18.48891, 15.66118, 12.24169,
    10.87285,
  10.39343, 10.14829, 10.36233, 10.64816, 10.92725, 11.04502, 10.95091,
    10.79418, 11.26044, 11.70811, 11.61377, 11.33595, 10.98827, 11.10115,
    11.69882, 12.05157, 11.15856, 10.52173, 10.80323, 14.98617, 16.51548,
    12.71474, 12.63737, 14.76434, 16.2927, 15.97144, 15.40558, 15.62723,
    15.60433, 11.94138,
  10.33427, 10.3314, 10.96429, 11.96908, 12.00569, 11.41168, 11.30326,
    11.10088, 10.88056, 11.01805, 10.93946, 12.185, 13.61234, 13.72145,
    13.01539, 18.56298, 23.97427, 17.56001, 13.46319, 15.86325, 14.65369,
    11.65092, 12.16819, 12.7647, 15.08933, 14.67026, 16.56723, 26.80258,
    23.69785, 11.56779,
  10.39082, 10.66148, 11.41311, 12.36442, 12.54419, 12.02116, 12.32348,
    13.54152, 13.77892, 13.72203, 14.31641, 14.12839, 13.30638, 13.17057,
    17.55482, 24.37145, 22.74159, 15.84457, 13.79245, 13.72504, 12.45121,
    11.64888, 12.07216, 14.00619, 15.42798, 13.13598, 21.35117, 35.33785,
    24.99834, 10.40502,
  10.5429, 10.83544, 11.69923, 12.54161, 12.44842, 14.2132, 15.99434,
    14.28667, 13.22465, 13.44038, 13.56019, 12.73877, 11.81467, 11.9377,
    14.46695, 16.55351, 15.22874, 13.69557, 12.64336, 12.42623, 11.92043,
    11.61843, 12.65695, 14.79265, 14.67589, 12.6951, 25.19753, 31.51875,
    16.49912, 10.63021,
  11.88853, 11.99065, 13.01695, 13.16238, 13.54156, 15.46598, 14.82689,
    13.15121, 13.25467, 13.49516, 13.00606, 12.18386, 11.75473, 14.86572,
    16.56967, 13.79489, 13.78994, 15.05033, 15.00949, 13.26401, 11.60707,
    12.55789, 15.97322, 16.95292, 14.2529, 14.18688, 20.97834, 20.5687,
    12.40945, 10.71963,
  13.951, 15.17551, 16.63804, 17.7301, 18.04126, 15.63674, 12.49699,
    12.33679, 12.27571, 11.81449, 13.01127, 16.29581, 17.77164, 17.67325,
    16.63725, 16.35498, 16.88233, 17.27368, 16.36812, 15.17644, 14.91043,
    15.68552, 16.98482, 15.81846, 19.79086, 28.15579, 23.01734, 13.55027,
    11.27228, 10.10328,
  22.99944, 26.14013, 23.59902, 19.3393, 18.68892, 17.72182, 14.84305,
    16.33346, 17.70404, 24.03396, 27.43751, 18.2345, 15.62649, 15.21667,
    14.64323, 15.51572, 16.66635, 16.54608, 15.46765, 15.34197, 17.4807,
    17.48368, 15.07943, 13.2728, 17.32508, 21.99756, 16.75942, 10.95934,
    10.38335, 9.92291,
  35.8845, 27.27371, 27.87415, 28.13479, 26.87782, 23.16182, 25.87331,
    24.0426, 19.53445, 24.31536, 24.4163, 14.00658, 14.79203, 15.78186,
    14.69065, 15.12347, 14.57662, 14.49757, 14.16273, 14.75565, 17.38829,
    16.54804, 12.89103, 15.62435, 17.73352, 12.9894, 10.3868, 10.62912,
    10.56291, 10.09032,
  42.29695, 38.54479, 53.60086, 58.45739, 58.17512, 49.6366, 36.46416,
    23.24138, 21.44454, 20.52771, 17.58671, 12.06376, 16.5268, 19.04899,
    15.73718, 15.08724, 15.01202, 14.4313, 14.05444, 16.33582, 17.96478,
    15.10601, 12.44068, 17.36093, 19.12753, 12.04595, 10.42606, 10.77809,
    11.04009, 10.38494,
  50.57007, 72.73684, 72.72933, 67.38799, 56.76711, 48.5619, 43.46455,
    37.11151, 29.86023, 25.88831, 30.62358, 30.34562, 34.1452, 34.36855,
    28.37224, 20.57184, 15.39067, 16.7078, 18.01681, 19.35383, 17.19886,
    16.17488, 17.97354, 15.70623, 13.21635, 10.99925, 10.51434, 10.41011,
    10.8204, 10.38732,
  37.25079, 44.99555, 42.9695, 40.07825, 33.8445, 38.01712, 53.88199,
    51.17146, 41.85104, 42.41781, 42.55604, 32.02047, 24.31392, 29.44359,
    31.29849, 19.57631, 18.59342, 18.4081, 20.26671, 21.83835, 19.79679,
    17.48891, 15.34839, 12.43731, 10.59395, 10.93876, 10.5492, 10.27598,
    10.33385, 10.12392,
  26.86124, 26.85961, 26.77055, 25.94688, 25.1416, 30.00592, 37.10056,
    34.6396, 31.64069, 31.76168, 29.07302, 21.41403, 16.4681, 20.68379,
    21.2338, 18.40444, 19.89806, 18.04805, 18.34337, 18.90914, 15.926,
    13.74283, 11.45565, 11.19835, 11.21868, 10.88189, 10.57647, 10.38733,
    10.26985, 10.04436,
  25.21275, 24.49185, 23.43132, 22.79538, 23.24267, 24.31181, 24.91587,
    24.47796, 23.98697, 22.66261, 18.54845, 17.81119, 20.08251, 18.68153,
    18.23234, 18.58454, 18.4533, 16.53418, 17.07324, 16.55655, 11.96756,
    11.85477, 11.70238, 11.51575, 11.18179, 10.94155, 10.55509, 10.21533,
    10.2006, 10.04643,
  22.67465, 22.00824, 21.08849, 21.33615, 21.80756, 22.72346, 23.26213,
    23.23009, 22.51206, 19.64875, 18.13718, 20.47026, 21.14187, 20.43598,
    22.06566, 20.53505, 17.05418, 14.65799, 16.53004, 15.70902, 11.73961,
    11.94339, 11.88793, 11.69036, 10.91953, 10.76153, 10.50496, 10.05774,
    10.04156, 9.968489,
  22.47942, 22.3857, 21.04144, 20.68253, 21.11089, 21.45457, 21.74043,
    21.47966, 19.9823, 18.0993, 19.58972, 20.30961, 17.35423, 18.0865,
    19.1153, 17.99022, 17.04719, 16.84834, 18.56282, 17.39399, 14.07591,
    12.75154, 11.93313, 11.65733, 10.74802, 10.50691, 10.40229, 10.06848,
    9.990678, 9.93623,
  22.96973, 23.0116, 21.49043, 20.33784, 20.57705, 20.59172, 20.50536, 20.08,
    19.06221, 19.94807, 20.88068, 17.6522, 15.29809, 15.36625, 15.14482,
    14.52769, 15.34037, 16.96714, 18.13484, 18.29436, 17.01344, 14.43828,
    12.02522, 11.63246, 10.96788, 10.50644, 10.35541, 10.11663, 9.998813,
    9.94091,
  22.70001, 22.90403, 21.42206, 20.24475, 20.14957, 20.13641, 20.01224,
    19.74306, 19.69911, 21.21319, 19.72518, 15.3004, 14.97185, 14.69771,
    13.8907, 13.21965, 13.43833, 14.20709, 14.98444, 15.39155, 15.79203,
    15.34417, 13.39207, 12.0785, 11.33904, 10.74659, 10.35396, 10.11537,
    10.01127, 9.946363,
  23.2083, 22.6624, 21.27445, 20.46099, 20.26727, 19.86889, 20.01977,
    20.00353, 20.74717, 21.04968, 17.54573, 14.0612, 14.05378, 13.74675,
    13.19277, 12.90079, 12.69636, 12.70693, 13.03073, 12.97027, 14.10068,
    14.43281, 13.3861, 13.67696, 12.69589, 11.17672, 10.4392, 10.1866,
    10.02298, 9.949555,
  23.20259, 22.78394, 21.13419, 20.29465, 20.79882, 21.23137, 21.4055,
    20.75418, 21.07512, 19.85284, 15.72047, 13.53963, 13.20148, 13.00147,
    12.61391, 12.85145, 12.88413, 12.27482, 12.0148, 11.91619, 13.16326,
    13.10512, 11.83103, 13.36511, 13.73817, 11.83403, 10.64198, 10.5823,
    10.24883, 9.964454,
  22.95872, 22.65321, 21.73806, 21.58597, 22.08318, 22.45248, 23.13712,
    23.06134, 22.81819, 19.42236, 14.97175, 13.8653, 13.61597, 13.74184,
    13.50245, 13.5713, 13.67371, 12.8375, 11.96971, 12.0312, 12.38308,
    12.07013, 11.49044, 11.88459, 12.86337, 13.13124, 11.93121, 10.88551,
    10.57809, 10.08823,
  23.16931, 23.96161, 22.14163, 21.76315, 22.56572, 22.80958, 22.68345,
    22.61991, 23.14637, 19.65124, 14.99148, 14.19086, 14.0263, 14.18353,
    14.21998, 14.17945, 13.65575, 13.15415, 12.49484, 12.01495, 11.96335,
    11.91075, 11.83377, 11.4247, 11.42389, 12.71892, 12.81758, 11.5789,
    11.41046, 10.51049,
  23.73083, 25.96017, 24.62002, 23.16934, 22.75264, 22.16563, 22.65174,
    23.39628, 22.27208, 18.81569, 15.54396, 14.70209, 14.57546, 14.23417,
    13.74034, 13.63789, 13.15405, 13.00049, 12.82709, 12.15035, 12.13618,
    12.22413, 11.62861, 11.15076, 11.12036, 11.78154, 13.09434, 12.32603,
    11.46944, 10.52118,
  24.97292, 27.47079, 25.14144, 23.0978, 22.18515, 21.18784, 22.69206,
    23.50071, 20.70084, 17.5171, 15.96968, 15.09612, 14.48126, 13.84861,
    13.39927, 13.18965, 12.86799, 12.85478, 12.7262, 12.09587, 12.16913,
    12.94149, 13.00018, 12.54927, 12.51372, 12.71365, 14.6268, 14.25075,
    11.4683, 10.06667,
  25.29396, 26.43889, 23.78029, 22.31037, 22.49757, 21.97279, 22.80472,
    22.11999, 18.8956, 17.06354, 15.83247, 14.73968, 13.84704, 13.54506,
    13.78985, 13.52925, 12.83395, 12.56918, 12.91229, 13.25599, 13.57466,
    13.6878, 13.41294, 13.03183, 13.19412, 13.28647, 14.00805, 15.65686,
    13.80476, 10.58285,
  23.36329, 22.45116, 22.1776, 23.14466, 23.94442, 24.46429, 23.72947,
    20.87359, 18.3115, 17.01051, 14.93426, 13.30114, 12.7077, 12.83008,
    13.41825, 13.63206, 13.46501, 13.66214, 13.50739, 13.18544, 13.24099,
    12.94983, 12.21488, 11.8408, 12.16132, 12.65124, 12.78995, 12.98568,
    13.3976, 11.15873,
  21.73005, 21.51497, 21.69353, 22.10427, 22.57112, 24.30005, 24.26828,
    20.63182, 17.73299, 16.62962, 15.16991, 14.34512, 14.2747, 14.25409,
    14.33308, 14.50752, 13.91031, 13.06818, 12.62497, 12.01701, 11.61986,
    11.54866, 11.32463, 11.22088, 11.34565, 11.9082, 12.05937, 11.42682,
    11.03214, 10.25514,
  12.78917, 12.80872, 12.83334, 12.8455, 12.84296, 12.83496, 12.82889,
    12.84442, 12.88342, 12.90454, 13.57033, 13.61794, 12.92332, 13.0761,
    13.16465, 12.92671, 12.86699, 12.88254, 12.86231, 13.24285, 13.46093,
    13.13139, 13.07063, 13.39299, 13.4403, 13.06881, 15.06053, 16.36433,
    14.40622, 13.38837,
  13.02129, 13.03055, 12.92825, 13.12277, 13.01029, 12.87804, 12.89448,
    12.92605, 12.99027, 13.11968, 13.54913, 13.93277, 14.03131, 13.57279,
    13.38143, 13.34061, 12.96223, 12.97236, 13.30275, 13.73883, 13.7193,
    13.16466, 13.03389, 13.48273, 16.36413, 16.66913, 16.34453, 19.19041,
    15.44804, 13.99114,
  13.02351, 13.02622, 12.98784, 13.069, 12.99581, 12.90495, 12.89429,
    12.96068, 13.05126, 13.12097, 13.1869, 13.51916, 13.79863, 14.04216,
    14.01086, 13.38903, 13.31628, 13.57944, 13.58352, 13.65241, 14.01983,
    14.80509, 15.52668, 14.90824, 19.24634, 21.87875, 18.30663, 18.9737,
    15.33911, 14.50568,
  12.96824, 12.95182, 13.10387, 13.21314, 13.38489, 13.73596, 13.71942,
    13.48631, 13.52051, 13.70335, 13.74458, 14.01914, 13.81527, 13.59259,
    14.24921, 14.87684, 14.39529, 13.58254, 13.49714, 13.43853, 15.4162,
    16.71532, 16.00024, 19.55072, 21.26617, 19.89269, 21.07435, 18.41049,
    15.16114, 13.89128,
  13.30158, 13.05548, 13.2659, 13.53492, 13.77979, 13.93248, 13.87854,
    13.67309, 14.08078, 14.51965, 14.45941, 14.2104, 13.86615, 13.94127,
    14.55813, 14.88817, 13.8567, 13.15989, 13.39772, 17.37938, 19.00906,
    15.46402, 15.28618, 17.47214, 18.92097, 18.44251, 18.08722, 18.40114,
    18.45539, 14.87076,
  13.23554, 13.18509, 13.80917, 14.80132, 14.84206, 14.26852, 14.18592,
    13.98642, 13.75215, 13.83482, 13.6655, 14.78081, 16.11801, 16.31452,
    15.52823, 20.48506, 25.70692, 19.92789, 15.94161, 18.51589, 17.47054,
    14.37797, 14.89234, 15.45045, 17.7225, 17.38061, 18.88461, 29.21794,
    26.83989, 14.54702,
  13.2194, 13.49211, 14.28662, 15.26358, 15.39888, 14.77625, 15.02114,
    16.1681, 16.307, 16.22787, 16.66862, 16.54791, 15.93207, 15.73112,
    19.82347, 26.76479, 25.65454, 18.70076, 16.54601, 16.51682, 15.20774,
    14.40839, 14.80136, 16.66202, 18.15377, 15.83975, 23.86756, 38.52033,
    28.58012, 13.33356,
  13.3638, 13.67103, 14.54777, 15.40308, 15.18121, 16.60411, 18.32362,
    16.93532, 15.98424, 16.13788, 16.20531, 15.35763, 14.41746, 14.42898,
    17.17705, 19.6097, 18.11089, 16.36227, 15.42914, 15.22503, 14.71612,
    14.4027, 15.34185, 17.46946, 17.46449, 15.32436, 28.30146, 35.20876,
    19.54909, 13.5182,
  14.51842, 14.60717, 15.63321, 15.79382, 16.00812, 17.99603, 17.56379,
    15.83056, 15.94142, 16.11417, 15.52519, 14.68871, 14.22167, 17.211,
    18.9375, 16.41532, 16.5045, 17.70799, 17.59168, 15.96566, 14.39115,
    15.24265, 18.49095, 19.48175, 16.86716, 16.68257, 23.95437, 23.80279,
    15.17716, 13.66157,
  16.16335, 17.26351, 18.86274, 20.06348, 20.31619, 18.00859, 15.06716,
    14.90471, 14.93578, 14.4033, 15.30926, 18.37195, 19.84583, 19.98337,
    19.17538, 18.83085, 19.33145, 19.67051, 18.90666, 17.93756, 17.65651,
    18.41397, 19.77128, 18.64426, 22.12289, 30.24247, 25.7637, 16.57665,
    14.28014, 13.06173,
  23.36133, 26.48208, 24.628, 20.79573, 20.51068, 19.60585, 16.85689,
    18.31347, 19.38197, 25.1221, 28.53052, 20.53197, 18.36868, 17.92408,
    17.26361, 18.15253, 19.33386, 19.23022, 18.18989, 18.2013, 20.37942,
    20.38833, 17.9796, 16.12886, 20.14175, 25.00576, 19.95747, 13.96604,
    13.3478, 12.86553,
  34.24454, 26.51449, 26.83948, 27.27323, 26.06452, 22.57365, 25.7733,
    24.70224, 20.58989, 25.55297, 26.20638, 16.5826, 17.32201, 18.35853,
    17.38814, 17.78826, 17.31108, 17.24216, 16.90394, 17.58469, 20.44074,
    19.63686, 15.82672, 18.47415, 20.69559, 16.08318, 13.37824, 13.54738,
    13.51599, 13.0448,
  39.67059, 33.43433, 44.49228, 50.35714, 50.57264, 44.58379, 34.20016,
    22.59993, 21.79595, 21.34746, 18.8167, 14.51471, 18.89065, 21.44189,
    18.45828, 17.76141, 17.7227, 17.1687, 16.78115, 19.25498, 21.15873,
    18.25054, 15.54015, 20.46779, 22.28109, 15.03707, 13.35018, 13.71639,
    13.99415, 13.339,
  44.87976, 63.87078, 66.1488, 66.22012, 61.94452, 51.63279, 37.34485,
    33.8362, 27.16185, 24.42734, 29.58648, 30.18349, 34.49191, 35.72536,
    30.83554, 23.26829, 18.19539, 19.55054, 20.93143, 22.46169, 20.36844,
    19.28075, 21.1646, 19.00751, 16.35688, 13.96979, 13.46539, 13.3771,
    13.80838, 13.36028,
  30.95862, 38.88078, 39.40468, 39.81472, 35.62217, 35.79253, 46.48671,
    45.9664, 36.76566, 38.16585, 39.76105, 31.71143, 26.36309, 31.58014,
    33.44142, 22.29103, 21.37064, 21.2671, 23.0433, 24.79937, 22.85369,
    20.59928, 18.53009, 15.5665, 13.61508, 13.98451, 13.56086, 13.26564,
    13.31246, 13.08695,
  20.47332, 20.61258, 21.39999, 21.10635, 19.51818, 23.71479, 31.48091,
    29.13142, 26.96523, 28.94216, 28.1832, 22.48901, 18.95911, 23.4001,
    23.82649, 21.19983, 22.85163, 21.06753, 21.19797, 21.91618, 19.07684,
    16.81625, 14.38873, 14.17892, 14.28084, 13.94397, 13.62348, 13.37572,
    13.2252, 12.98573,
  18.85502, 18.17002, 17.41496, 16.62495, 16.62934, 17.77886, 18.76681,
    18.52006, 19.13462, 19.96218, 18.15238, 19.1406, 22.27039, 21.29872,
    21.2145, 21.5892, 21.65124, 19.66008, 20.0546, 19.73187, 15.10299,
    14.9327, 14.6899, 14.50533, 14.16016, 13.96514, 13.56944, 13.19156,
    13.14726, 12.98063,
  16.417, 15.62372, 14.73879, 14.86269, 15.33568, 16.18831, 16.86909,
    17.36757, 17.64142, 16.75122, 17.29879, 21.48913, 23.60435, 23.30862,
    25.19274, 23.73093, 20.29646, 17.72987, 19.52408, 18.78377, 14.75188,
    14.95, 14.88792, 14.63808, 13.86226, 13.728, 13.48607, 13.01716,
    12.98723, 12.90792,
  16.18363, 15.82285, 14.46691, 14.06768, 14.52555, 14.94007, 15.28244,
    15.42429, 15.03523, 15.02062, 18.62682, 21.42544, 19.95808, 21.19287,
    22.37219, 21.1988, 20.16006, 19.58956, 21.30661, 20.32755, 17.04906,
    15.69919, 14.88627, 14.6067, 13.70027, 13.44162, 13.3568, 13.0286,
    12.93411, 12.86971,
  16.56902, 16.32918, 14.85329, 13.75025, 13.97287, 13.97357, 13.92396,
    13.87662, 13.96739, 16.7469, 20.00761, 18.96857, 17.88773, 18.38704,
    18.26476, 17.64457, 18.352, 19.81987, 20.99285, 21.32095, 19.91825,
    17.28828, 14.96117, 14.60054, 13.93303, 13.43854, 13.29835, 13.06458,
    12.93724, 12.8778,
  16.16757, 16.15086, 14.78996, 13.6117, 13.52871, 13.4805, 13.35054,
    13.4469, 14.5566, 18.10775, 19.05717, 16.70177, 17.60553, 17.73604,
    16.9209, 16.21232, 16.391, 17.16089, 17.97885, 18.42319, 18.90172,
    18.36665, 16.24424, 15.0544, 14.29578, 13.67235, 13.29486, 13.05202,
    12.94646, 12.88015,
  16.67175, 15.82902, 14.59023, 13.77806, 13.5785, 13.15657, 13.33154,
    13.74577, 15.71597, 18.20127, 17.08892, 15.40326, 16.58756, 16.71123,
    16.19719, 15.85345, 15.62854, 15.64828, 16.03497, 16.03557, 17.19718,
    17.44993, 16.36465, 16.59921, 15.4794, 14.01597, 13.34073, 13.10866,
    12.95436, 12.87703,
  16.74592, 15.88925, 14.33916, 13.57718, 14.06711, 14.48967, 14.79716,
    14.65954, 16.14138, 16.96914, 15.16622, 14.77256, 15.62048, 15.87941,
    15.59019, 15.80666, 15.77524, 15.17482, 14.98086, 14.96949, 16.17969,
    16.05014, 14.81474, 16.23063, 16.49956, 14.68712, 13.51762, 13.47711,
    13.1881, 12.90142,
  16.42468, 15.79245, 14.90429, 14.77413, 15.41351, 15.9101, 16.83967,
    17.31287, 17.93958, 16.24209, 14.17702, 14.97198, 15.86757, 16.49808,
    16.34176, 16.37637, 16.49083, 15.66399, 14.85202, 14.95756, 15.28342,
    14.94393, 14.3636, 14.72157, 15.7164, 15.96016, 14.73341, 13.76646,
    13.51607, 13.02626,
  16.46516, 16.589, 15.22238, 15.13835, 16.21403, 16.75294, 16.80052,
    16.90724, 18.07185, 16.32093, 14.01168, 15.2226, 16.271, 16.88678,
    16.97689, 16.91721, 16.48929, 16.00088, 15.34452, 14.90638, 14.79974,
    14.72871, 14.68778, 14.30594, 14.35641, 15.69629, 15.77513, 14.51142,
    14.31604, 13.43392,
  16.91057, 18.29954, 17.5778, 16.69168, 16.66898, 16.5198, 16.92528,
    17.50689, 16.94118, 15.41791, 14.44537, 15.69622, 16.83256, 16.91238,
    16.5083, 16.43366, 16.00516, 15.8416, 15.6754, 15.05645, 14.97725,
    15.09154, 14.53246, 14.05813, 14.0701, 14.79523, 16.10491, 15.29146,
    14.365, 13.42859,
  18.19289, 19.92904, 18.47491, 16.98127, 16.21386, 15.49411, 17.1434,
    17.86576, 15.41898, 14.12776, 14.95095, 16.16935, 16.83962, 16.61626,
    16.20107, 15.97727, 15.70122, 15.70295, 15.56712, 14.99373, 15.04475,
    15.87246, 15.93569, 15.46308, 15.51414, 15.7712, 17.6914, 17.27267,
    14.36573, 12.95604,
  19.01674, 19.79693, 17.45785, 16.27651, 16.35645, 15.86817, 16.80698,
    16.19108, 13.63884, 13.67029, 14.95757, 16.03728, 16.38013, 16.34047,
    16.51992, 16.27252, 15.64273, 15.41354, 15.78715, 16.20293, 16.48191,
    16.5917, 16.35446, 16.00598, 16.25575, 16.37738, 17.06607, 18.69255,
    16.76247, 13.49428,
  17.7023, 16.52143, 16.19569, 17.21194, 17.72878, 17.77175, 17.08825,
    14.5432, 12.96968, 13.66896, 14.22493, 14.78717, 15.2843, 15.67803,
    16.28284, 16.52583, 16.40384, 16.53979, 16.4349, 16.23289, 16.26031,
    15.90784, 15.17203, 14.83616, 15.17882, 15.66685, 15.77121, 16.03434,
    16.3919, 14.08812,
  16.86465, 16.2781, 16.41886, 16.90707, 17.10136, 18.22032, 17.98811,
    14.71041, 12.93272, 13.84166, 14.80377, 15.94896, 16.80207, 16.99485,
    17.12322, 17.37951, 16.8438, 16.03982, 15.65465, 15.04788, 14.63107,
    14.54724, 14.30955, 14.20365, 14.324, 14.88189, 15.03812, 14.41132,
    14.00687, 13.20086,
  12.62708, 12.64621, 12.67685, 12.69138, 12.68927, 12.6798, 12.6714,
    12.68499, 12.70603, 12.7223, 13.37487, 13.47644, 12.75546, 12.90355,
    13.0049, 12.76504, 12.72415, 12.74261, 12.71734, 13.1168, 13.35536,
    12.99885, 12.92111, 13.22789, 13.27594, 12.86579, 14.88832, 16.49756,
    14.45651, 13.35722,
  12.87941, 12.90946, 12.76483, 12.98439, 12.87124, 12.72934, 12.74547,
    12.76322, 12.80906, 12.93648, 13.42423, 13.85128, 13.90981, 13.47587,
    13.25785, 13.23883, 12.83883, 12.8373, 13.1956, 13.71877, 13.71195,
    13.07641, 12.84174, 13.27681, 16.1154, 16.76604, 16.35981, 19.81368,
    15.71202, 14.09937,
  12.9045, 12.90985, 12.84373, 12.94707, 12.86439, 12.743, 12.72157,
    12.79227, 12.88462, 12.96231, 13.03725, 13.42358, 13.77862, 14.00311,
    13.9736, 13.3004, 13.1747, 13.50426, 13.5541, 13.63043, 13.93817,
    14.66679, 15.3334, 14.62973, 19.1131, 22.75343, 18.59747, 19.69809,
    15.57344, 14.65197,
  12.83683, 12.80545, 12.94506, 13.03774, 13.21015, 13.58239, 13.59237,
    13.36595, 13.35798, 13.53529, 13.62648, 13.92681, 13.75479, 13.53165,
    14.22143, 14.91401, 14.50683, 13.56848, 13.38174, 13.20517, 15.15266,
    16.66731, 15.79451, 19.54004, 21.99911, 20.3253, 21.77437, 19.10409,
    15.37748, 13.92778,
  13.18158, 12.88897, 13.06569, 13.32756, 13.65209, 13.89367, 13.82001,
    13.56282, 13.95867, 14.49641, 14.49099, 14.18032, 13.72862, 13.82719,
    14.59243, 15.04971, 13.91852, 12.94407, 13.08473, 17.01136, 19.11321,
    15.39993, 15.07851, 17.57262, 19.34805, 18.79935, 18.69414, 18.9418,
    18.86649, 14.93272,
  13.0993, 12.97588, 13.54622, 14.56169, 14.79364, 14.29089, 14.09107,
    13.85745, 13.6846, 13.79974, 13.59186, 14.63389, 16.0713, 16.30068,
    15.62218, 20.40916, 26.15982, 20.29004, 15.61984, 18.43526, 17.69112,
    14.23383, 14.78121, 15.45919, 17.93469, 17.88688, 18.77503, 29.39244,
    27.76051, 14.68295,
  13.00241, 13.22621, 14.0384, 15.10772, 15.39303, 14.79863, 14.88092,
    16.08323, 16.14112, 15.97473, 16.52983, 16.58746, 16.0407, 15.73791,
    19.83544, 27.54679, 26.92712, 19.14058, 16.47079, 16.5468, 15.20082,
    14.32567, 14.76605, 16.75619, 18.44079, 16.02268, 23.81396, 39.92284,
    30.33352, 13.32441,
  13.12972, 13.43933, 14.32403, 15.22715, 15.08272, 16.44877, 18.31614,
    17.02541, 15.85561, 16.0518, 16.32866, 15.46644, 14.28775, 14.19284,
    17.22942, 20.30041, 18.57248, 16.40424, 15.36724, 15.20992, 14.71407,
    14.37298, 15.35771, 17.64667, 17.71021, 15.31021, 28.8374, 37.49133,
    20.31687, 13.48216,
  14.21543, 14.31571, 15.27118, 15.49622, 15.7507, 18.09435, 17.90237,
    15.80506, 15.79359, 16.08363, 15.53326, 14.51987, 13.82741, 16.90118,
    19.10393, 16.52452, 16.59036, 18.00594, 17.81265, 16.07716, 14.34359,
    15.27285, 18.68173, 19.88286, 17.03568, 16.66318, 24.46542, 24.92053,
    15.09387, 13.61522,
  15.96754, 16.97586, 18.63961, 20.05894, 20.32059, 18.22852, 15.16587,
    14.84091, 14.83914, 14.24489, 14.96607, 18.16698, 19.82558, 20.14605,
    19.43698, 18.99258, 19.56826, 20.14821, 19.44726, 18.28095, 17.87004,
    18.70958, 20.20962, 19.0514, 22.25373, 30.59178, 26.39936, 16.84609,
    14.24281, 12.93261,
  22.23582, 25.78115, 24.78527, 21.06498, 20.76796, 20.02511, 17.11235,
    18.48059, 19.27419, 24.67984, 28.78879, 20.8534, 18.61309, 18.1414,
    17.36997, 18.36435, 19.8168, 19.79424, 18.69612, 18.59342, 20.85851,
    20.87132, 18.29795, 16.24808, 20.44127, 25.82092, 20.7131, 14.00865,
    13.21804, 12.70436,
  35.56506, 28.46991, 26.88039, 27.22961, 26.13877, 22.50794, 25.73116,
    25.20738, 20.92013, 25.77527, 27.01253, 16.67789, 17.25429, 18.52262,
    17.6279, 18.13552, 17.7129, 17.61941, 17.20665, 17.88875, 20.87699,
    20.02442, 15.91434, 18.49, 21.20036, 16.60867, 13.43941, 13.41195,
    13.38051, 12.89889,
  49.94715, 38.9021, 42.54939, 50.02816, 50.40609, 45.51487, 36.20273,
    23.3727, 22.56394, 22.06238, 19.55315, 14.31981, 18.80934, 21.82224,
    18.87783, 18.04956, 18.06002, 17.49091, 16.97732, 19.61206, 21.73704,
    18.4678, 15.60028, 20.79153, 23.20992, 15.29778, 13.24469, 13.59924,
    13.91197, 13.26432,
  51.38953, 65.67749, 65.72362, 68.29703, 63.84121, 54.30443, 40.39191,
    36.08812, 29.30043, 24.83642, 30.17068, 30.65394, 35.05098, 35.51514,
    30.48309, 23.79615, 18.43107, 19.93235, 21.58556, 23.26217, 20.91948,
    19.59916, 21.92628, 19.65376, 16.87123, 13.98601, 13.36654, 13.27865,
    13.75016, 13.29457,
  33.80087, 40.73561, 41.62389, 43.75278, 39.90739, 38.87816, 48.68777,
    48.53829, 37.91682, 38.23363, 40.44706, 33.25999, 27.10855, 31.64573,
    33.86555, 22.68794, 21.7459, 21.7872, 23.82301, 25.89286, 23.80184,
    21.46282, 19.37463, 15.98485, 13.54975, 13.90551, 13.471, 13.18277,
    13.22962, 12.9788,
  22.79552, 23.13309, 24.575, 24.8079, 23.06382, 26.84112, 34.50198,
    31.51958, 28.59507, 30.44005, 29.8406, 23.91103, 19.73164, 24.31358,
    24.55687, 21.60756, 23.45528, 21.68908, 21.85913, 22.86751, 19.86849,
    17.44253, 14.6375, 14.24609, 14.25383, 13.89341, 13.55401, 13.28913,
    13.11482, 12.85528,
  21.51112, 21.09969, 20.5687, 19.62962, 19.37435, 20.681, 21.93589,
    21.40756, 21.75781, 22.47572, 19.99397, 20.21083, 23.21282, 22.07635,
    21.86782, 22.10487, 22.2866, 20.23927, 20.68474, 20.58305, 15.37488,
    15.09451, 14.71321, 14.51817, 14.14724, 13.92377, 13.5057, 13.08555,
    13.02048, 12.84431,
  19.14228, 18.56346, 17.5542, 17.59363, 18.07622, 19.00818, 19.7954,
    20.32068, 20.41895, 18.9789, 18.616, 22.51441, 24.52099, 23.85928,
    26.34771, 24.68363, 20.95437, 18.07319, 20.1262, 19.59318, 14.82657,
    14.97132, 14.84953, 14.63195, 13.79759, 13.65759, 13.42165, 12.88562,
    12.85068, 12.7647,
  18.99144, 18.68409, 17.21196, 16.79555, 17.26354, 17.76194, 18.26144,
    18.43627, 17.81873, 17.04745, 19.91913, 22.42165, 20.4599, 21.69835,
    23.52181, 22.34109, 21.00249, 19.97792, 21.85908, 20.76675, 16.93454,
    15.65317, 14.85949, 14.57752, 13.60836, 13.35133, 13.27836, 12.89934,
    12.79386, 12.71973,
  19.43764, 19.20579, 17.65028, 16.48165, 16.75052, 16.8417, 16.91831,
    16.86067, 16.57425, 18.7459, 21.56769, 19.93815, 18.27827, 18.87524,
    19.05585, 18.52434, 19.26149, 20.45129, 21.26858, 21.53053, 19.96826,
    17.42172, 14.94338, 14.55444, 13.86936, 13.35107, 13.20194, 12.93896,
    12.79215, 12.72698,
  18.93662, 18.97141, 17.6144, 16.42434, 16.38975, 16.44549, 16.34481,
    16.31376, 17.12617, 20.36254, 20.88384, 17.64769, 18.12983, 18.256,
    17.50025, 16.70319, 16.83003, 17.37115, 18.01996, 18.66554, 19.27946,
    18.73633, 16.27572, 15.09683, 14.32366, 13.62727, 13.18661, 12.91751,
    12.79892, 12.73471,
  19.41562, 18.63685, 17.47687, 16.70401, 16.53733, 16.10019, 16.25217,
    16.61226, 18.41674, 20.68159, 19.01295, 16.44581, 17.27253, 17.23565,
    16.55638, 16.02625, 15.67869, 15.61885, 16.12078, 16.2199, 17.47081,
    17.8847, 16.52734, 16.82487, 15.65056, 14.01297, 13.21889, 12.98207,
    12.8025, 12.72646,
  19.57633, 18.7926, 17.32597, 16.55247, 17.02552, 17.39899, 17.70667,
    17.59349, 19.07227, 19.70722, 17.1369, 15.92273, 16.27372, 16.2145,
    15.71314, 15.82298, 15.80436, 15.24415, 15.07669, 15.02777, 16.38608,
    16.4452, 14.95067, 16.51301, 16.79838, 14.79419, 13.43274, 13.37244,
    13.05763, 12.75433,
  19.43045, 18.83343, 17.89828, 17.72038, 18.37343, 18.91808, 20.00882,
    20.68127, 21.42506, 19.25191, 16.14131, 16.0873, 16.30711, 16.59985,
    16.34568, 16.39741, 16.6354, 15.81511, 14.8856, 15.03606, 15.55448,
    15.20922, 14.44611, 14.86208, 15.93878, 16.11272, 14.72846, 13.68399,
    13.41834, 12.90077,
  19.39849, 19.38251, 18.10813, 18.0688, 19.23836, 20.10776, 20.50593,
    20.74215, 21.90124, 19.53158, 15.82986, 16.19572, 16.65006, 17.01782,
    17.04304, 17.09342, 16.73542, 16.17554, 15.41413, 15.03272, 15.01553,
    14.87868, 14.78728, 14.37201, 14.40547, 15.80006, 15.89303, 14.52249,
    14.27433, 13.37437,
  19.76722, 20.82965, 20.35674, 19.76972, 19.96191, 20.20906, 20.79391,
    21.53478, 20.72355, 18.39981, 16.05856, 16.52554, 17.25736, 17.17895,
    16.67787, 16.60532, 16.16997, 15.94073, 15.75704, 15.19889, 15.15681,
    15.22731, 14.59257, 14.0324, 14.00092, 14.8032, 16.21783, 15.38821,
    14.33764, 13.38801,
  20.98253, 22.33996, 21.4908, 20.4873, 19.79542, 19.16014, 20.94058,
    21.7768, 18.85381, 16.63881, 16.47235, 16.99344, 17.31112, 16.90817,
    16.3267, 16.04825, 15.79556, 15.80917, 15.68061, 15.11274, 15.19253,
    16.07167, 16.09517, 15.47015, 15.42778, 15.68158, 17.73102, 17.39776,
    14.34671, 12.8707,
  22.18295, 22.77282, 20.5746, 19.95, 20.03466, 19.49278, 20.52014, 19.78018,
    16.64782, 15.93596, 16.43521, 16.84941, 16.78083, 16.51678, 16.58722,
    16.31549, 15.68993, 15.49283, 15.90604, 16.35991, 16.70829, 16.88133,
    16.54667, 16.05218, 16.20287, 16.3688, 17.177, 18.90581, 16.99762,
    13.47589,
  21.15707, 19.93586, 19.5983, 20.87456, 21.4378, 21.44323, 20.7761,
    17.94663, 15.86442, 15.99197, 15.74788, 15.54215, 15.52294, 15.71878,
    16.30679, 16.53454, 16.41532, 16.59827, 16.61448, 16.50616, 16.51694,
    16.08373, 15.23536, 14.80437, 15.13961, 15.67599, 15.84095, 16.20745,
    16.65745, 14.1816,
  20.12018, 19.54296, 19.74644, 20.23116, 20.50433, 21.78526, 21.48852,
    17.92413, 15.69228, 16.04352, 16.18139, 16.55808, 16.96132, 17.08455,
    17.20331, 17.42581, 16.92653, 16.10224, 15.76516, 15.18209, 14.68554,
    14.56357, 14.29422, 14.14202, 14.25251, 14.81994, 15.02712, 14.39979,
    14.01059, 13.14597,
  16.11749, 16.13822, 16.15806, 16.17335, 16.17391, 16.16201, 16.16579,
    16.18361, 16.19895, 16.21517, 16.86402, 17.01341, 16.26208, 16.42765,
    16.57563, 16.31036, 16.24946, 16.25582, 16.22131, 16.63954, 16.91857,
    16.5376, 16.45852, 16.7977, 16.81847, 16.36753, 18.44728, 20.24484,
    18.18783, 17.02018,
  16.366, 16.40318, 16.24761, 16.49257, 16.3786, 16.22542, 16.2422, 16.26469,
    16.30325, 16.44308, 17.00703, 17.50034, 17.56402, 17.12688, 16.88948,
    16.87056, 16.38077, 16.35867, 16.75673, 17.38904, 17.43637, 16.68885,
    16.36623, 16.88667, 19.62068, 20.3112, 20.32699, 24.44983, 19.82338,
    17.90672,
  16.43318, 16.44575, 16.36536, 16.49322, 16.3831, 16.24853, 16.21954,
    16.27272, 16.39276, 16.51254, 16.62213, 17.07479, 17.51184, 17.69476,
    17.64119, 16.93515, 16.73245, 17.12227, 17.23479, 17.34083, 17.63887,
    18.38293, 19.06439, 18.29638, 22.93021, 27.1495, 22.98241, 24.62631,
    19.6228, 18.49617,
  16.34716, 16.33411, 16.48262, 16.57924, 16.75752, 17.17826, 17.18957,
    16.91491, 16.90974, 17.09459, 17.213, 17.59016, 17.4235, 17.13629,
    17.9089, 18.66245, 18.2775, 17.26734, 17.01531, 16.72486, 18.85898,
    20.70939, 19.62657, 23.57756, 26.54274, 25.022, 26.9129, 23.77997,
    19.32889, 17.72364,
  16.7496, 16.43073, 16.60507, 16.86546, 17.24309, 17.60021, 17.52641,
    17.18116, 17.57554, 18.21921, 18.31831, 17.9307, 17.34031, 17.41596,
    18.25091, 18.88979, 17.6894, 16.42077, 16.4959, 20.68483, 23.37669,
    19.24532, 18.73524, 21.74659, 23.95021, 23.29301, 23.40738, 23.41853,
    23.17447, 18.78842,
  16.70088, 16.49885, 17.1126, 18.19005, 18.46321, 17.95261, 17.70354,
    17.4745, 17.3271, 17.49868, 17.2549, 18.27774, 19.93534, 20.19098,
    19.43668, 23.88425, 29.88924, 24.18564, 19.34703, 22.68363, 22.00827,
    17.7398, 18.42554, 19.35243, 22.22518, 22.36433, 22.75031, 34.47275,
    33.56405, 18.64317,
  16.52704, 16.74455, 17.71415, 18.93975, 19.23987, 18.54127, 18.45451,
    19.80549, 19.97214, 19.78928, 20.36367, 20.50854, 20.02499, 19.63703,
    23.79338, 32.24253, 31.98521, 23.51374, 20.56618, 20.70956, 19.01212,
    17.91568, 18.50943, 20.8048, 22.80708, 20.14597, 27.83093, 46.55414,
    37.58681, 17.11127,
  16.65991, 17.01244, 18.05785, 19.09821, 18.90786, 20.25448, 22.35182,
    21.14377, 19.84717, 20.07147, 20.48743, 19.50484, 17.9742, 17.75704,
    21.27083, 25.11684, 23.08091, 20.47822, 19.26808, 19.08135, 18.46656,
    18.08368, 19.24136, 21.8793, 21.96351, 19.08067, 34.00622, 45.51169,
    25.92302, 17.2037,
  17.81439, 17.99852, 19.03823, 19.25245, 19.51188, 22.41893, 22.44433,
    19.82795, 19.70026, 20.10773, 19.55288, 18.27622, 17.3297, 20.55301,
    23.21276, 20.51807, 20.56803, 22.29534, 21.98088, 20.05634, 18.093,
    19.13357, 22.96153, 24.34991, 20.96918, 20.39261, 29.97726, 31.47658,
    19.11345, 17.39336,
  19.92537, 20.7357, 22.5752, 24.48877, 24.75769, 22.58398, 19.14556,
    18.69896, 18.78073, 18.12724, 18.71641, 22.10448, 23.7597, 24.29302,
    23.74734, 23.13354, 23.78698, 24.6144, 23.97021, 22.41105, 21.82646,
    22.93056, 24.82302, 23.4596, 26.24083, 35.54901, 32.07802, 21.55425,
    18.23981, 16.58508,
  25.54593, 29.76829, 29.27406, 25.17808, 25.13058, 24.5323, 21.42686,
    22.7069, 23.64084, 28.7923, 33.34508, 25.36427, 22.87101, 22.25097,
    21.22982, 22.50951, 24.31976, 24.27793, 23.00363, 22.7187, 25.31507,
    25.57701, 22.75023, 20.14698, 24.8767, 31.7868, 26.35137, 18.05688,
    16.93853, 16.24175,
  40.27147, 33.0138, 30.51478, 30.34872, 29.81786, 25.28415, 29.2431,
    29.97239, 25.54478, 30.79416, 32.48262, 20.71837, 20.95301, 22.26253,
    21.54153, 22.25699, 21.924, 21.80626, 21.26585, 21.98384, 25.47239,
    24.68569, 19.97433, 22.4714, 25.94046, 21.30151, 17.43253, 17.13433,
    17.0498, 16.45369,
  53.63425, 39.56782, 43.24854, 50.3175, 52.87835, 50.68343, 43.40244,
    27.88971, 28.14568, 27.43359, 24.0458, 17.74794, 22.52851, 25.76832,
    22.98783, 22.15269, 22.29188, 21.52118, 20.82547, 23.73111, 26.40379,
    22.75008, 19.49079, 25.50344, 28.93849, 19.66392, 16.92119, 17.32755,
    17.6542, 16.89801,
  54.7649, 59.24383, 59.70531, 64.96871, 65.28175, 61.24615, 47.16397,
    41.47412, 35.26495, 28.86374, 34.23058, 33.90625, 39.39433, 40.28901,
    35.20805, 28.12518, 22.71125, 24.37719, 26.0482, 27.96305, 25.59867,
    23.68498, 26.77584, 25.12589, 21.91758, 17.88678, 17.01579, 16.95969,
    17.51342, 16.97009,
  37.17351, 41.35193, 45.28957, 52.01309, 53.85854, 49.62459, 52.21927,
    53.46939, 40.89381, 40.66055, 43.74589, 37.93142, 32.09318, 36.9822,
    39.08258, 27.46235, 26.33662, 26.57063, 28.80355, 30.78213, 28.10354,
    26.08928, 24.70594, 20.84063, 17.36397, 17.69847, 17.14197, 16.81259,
    16.89099, 16.58646,
  25.79149, 28.45068, 33.16588, 35.70869, 33.91014, 33.15454, 37.74429,
    34.55781, 30.71533, 33.35944, 33.42782, 27.86697, 23.44263, 29.0161,
    29.41062, 26.06128, 28.30495, 26.39818, 26.55203, 27.78707, 24.60628,
    22.16402, 18.90471, 18.09177, 17.98418, 17.65389, 17.2307, 16.94033,
    16.73721, 16.42038,
  23.778, 24.52866, 24.86008, 23.55144, 21.88329, 22.56311, 24.12494,
    23.21042, 23.68205, 25.02357, 22.58763, 22.79329, 26.55088, 26.05205,
    26.21493, 26.5569, 26.97146, 24.77389, 25.26406, 25.66798, 19.84608,
    19.25398, 18.53343, 18.21083, 17.85977, 17.70258, 17.22219, 16.71874,
    16.6418, 16.41599,
  20.59414, 20.1392, 18.88256, 18.35329, 18.56781, 19.80018, 20.73576,
    21.36077, 21.76172, 20.38082, 19.95329, 24.76606, 27.97837, 27.67334,
    31.25624, 29.51403, 25.47764, 22.44807, 25.01889, 24.79859, 18.9846,
    18.88677, 18.59066, 18.33723, 17.48796, 17.41964, 17.15711, 16.49394,
    16.42701, 16.31437,
  19.96415, 19.4656, 17.63227, 17.05805, 17.55771, 18.10876, 18.6948,
    18.99073, 18.43779, 17.47895, 20.91771, 24.65109, 23.40981, 25.62439,
    28.56535, 27.18162, 25.57293, 24.42188, 26.94674, 25.64537, 20.86338,
    19.46465, 18.64648, 18.34997, 17.29243, 17.00367, 16.93092, 16.48974,
    16.35033, 16.26209,
  20.24431, 19.63159, 17.78724, 16.43307, 16.75733, 16.92323, 17.12311,
    17.11848, 16.62694, 18.91613, 22.62238, 21.80589, 20.80276, 22.51932,
    23.46203, 23.00871, 23.91542, 25.35727, 26.28388, 26.32233, 24.24386,
    21.46574, 18.78735, 18.36763, 17.56663, 16.97742, 16.8191, 16.51882,
    16.33779, 16.26408,
  19.45691, 19.16543, 17.66134, 16.3563, 16.38068, 16.54478, 16.4591,
    16.25879, 16.97553, 20.72827, 22.04616, 19.26265, 20.79746, 21.89764,
    21.66247, 21.09142, 21.35461, 21.97016, 22.4653, 23.16582, 23.91065,
    23.15682, 20.18087, 18.93676, 18.02128, 17.28214, 16.80468, 16.49154,
    16.33802, 16.26088,
  19.89531, 18.76542, 17.52106, 16.73577, 16.62289, 16.16092, 16.19377,
    16.39373, 18.42909, 21.3146, 20.08795, 18.04112, 20.00175, 20.8992,
    20.76173, 20.36894, 19.93897, 19.74449, 20.30075, 20.43731, 21.85256,
    22.42696, 20.67518, 20.92064, 19.50407, 17.73028, 16.8252, 16.54778,
    16.34832, 16.26553,
  20.14415, 18.97014, 17.41529, 16.63879, 17.16484, 17.40191, 17.59907,
    17.47868, 19.41249, 20.63767, 18.1757, 17.56616, 19.01411, 19.80383,
    19.76043, 20.045, 19.95819, 19.26491, 19.11463, 19.01352, 20.549,
    20.72927, 18.99362, 20.85639, 21.01237, 18.61742, 17.04561, 17.01331,
    16.64346, 16.29005,
  19.99315, 19.0999, 18.12443, 17.8317, 18.45726, 18.94932, 20.17092,
    21.13707, 22.23857, 20.17666, 17.06966, 17.79802, 19.06046, 20.13375,
    20.27122, 20.47108, 20.76877, 19.91717, 18.82634, 18.85792, 19.54497,
    19.21856, 18.28991, 18.94046, 20.16076, 20.06294, 18.44556, 17.42298,
    17.08825, 16.45938,
  19.99472, 19.75053, 18.3519, 18.12545, 19.28256, 20.32595, 21.0679,
    21.68307, 23.1025, 20.56748, 16.81756, 18.04077, 19.37961, 20.52575,
    21.02269, 21.25865, 21.00453, 20.33657, 19.33992, 18.89033, 18.8867,
    18.72674, 18.6553, 18.207, 18.25784, 19.78446, 19.79771, 18.31082,
    18.04544, 17.01289,
  20.29197, 21.14407, 20.41638, 19.6851, 20.03878, 20.67922, 21.6587,
    22.70114, 21.86332, 19.44691, 17.06373, 18.32086, 19.92802, 20.67069,
    20.66425, 20.82336, 20.35991, 19.93739, 19.66859, 19.068, 19.05326,
    19.187, 18.48269, 17.75127, 17.6417, 18.58395, 20.10508, 19.23464,
    18.14241, 17.06119,
  21.40081, 22.54774, 21.7647, 20.68332, 20.12198, 19.74182, 22.12569,
    23.35271, 19.90323, 17.41398, 17.42607, 18.72458, 20.08742, 20.55109,
    20.38204, 20.13657, 19.73009, 19.65826, 19.54659, 18.98372, 19.14144,
    20.11666, 20.06124, 19.24333, 19.09716, 19.38861, 21.59666, 21.3314,
    18.07684, 16.4386,
  22.76628, 23.42571, 20.92635, 20.33335, 20.61843, 20.3801, 21.88801,
    21.25467, 17.38755, 16.4349, 17.31767, 18.62247, 19.62983, 20.19839,
    20.67505, 20.38737, 19.58698, 19.32856, 19.77771, 20.25695, 20.76293,
    21.10354, 20.70594, 20.04016, 20.04603, 20.24772, 21.21322, 23.10529,
    21.02811, 17.10305,
  21.78013, 20.45009, 20.18211, 22.00187, 22.72947, 22.73656, 22.16709,
    18.9732, 16.31507, 16.44481, 16.61654, 17.30764, 18.30897, 19.31739,
    20.4039, 20.668, 20.40021, 20.56393, 20.60922, 20.56232, 20.70398,
    20.25561, 19.21939, 18.64014, 18.99135, 19.61882, 19.83908, 20.44926,
    20.96936, 18.00691,
  20.91902, 20.3068, 20.96198, 21.90903, 22.11938, 23.39866, 22.96061,
    18.78385, 16.1699, 16.67909, 17.24421, 18.42033, 19.73088, 20.58865,
    21.24463, 21.65616, 21.07547, 20.21834, 19.83403, 19.09726, 18.5613,
    18.422, 18.06238, 17.86621, 18.02722, 18.699, 18.98419, 18.31405,
    17.95113, 16.85873,
  18.3728, 18.42345, 18.43662, 18.44517, 18.44161, 18.43993, 18.44011,
    18.46194, 18.478, 18.50613, 19.26756, 19.50903, 18.56127, 18.71857,
    18.88769, 18.56996, 18.49939, 18.52536, 18.51211, 18.99897, 19.39241,
    18.94682, 18.86769, 19.26106, 19.27766, 18.77813, 21.08584, 23.57801,
    21.0126, 19.62972,
  18.621, 18.72345, 18.52178, 18.80324, 18.66011, 18.48688, 18.51442,
    18.53153, 18.58537, 18.77884, 19.39267, 19.91937, 19.98964, 19.50217,
    19.15032, 19.19408, 18.65164, 18.63911, 19.14922, 19.9094, 19.91134,
    19.05338, 18.70188, 19.43005, 22.66469, 24.22407, 23.78901, 29.20087,
    22.96292, 20.7114,
  18.71304, 18.74632, 18.65299, 18.78045, 18.64508, 18.50124, 18.4804,
    18.56532, 18.69314, 18.82692, 18.96009, 19.41128, 19.87443, 20.09865,
    20.0552, 19.24687, 19.05912, 19.59453, 19.74866, 19.84708, 20.1688,
    21.12118, 21.91952, 21.38966, 26.45951, 32.13673, 27.36755, 29.39963,
    22.64771, 21.39299,
  18.62034, 18.60151, 18.77174, 18.90207, 19.10354, 19.6006, 19.60991,
    19.27948, 19.24778, 19.41196, 19.57746, 20.02785, 19.88294, 19.48291,
    20.41288, 21.41254, 21.13349, 19.85313, 19.42839, 19.13895, 21.61426,
    23.95523, 22.6875, 27.24678, 30.95996, 29.04649, 32.25948, 27.94088,
    22.32822, 20.39021,
  19.10141, 18.68095, 18.89916, 19.2097, 19.65497, 20.0462, 19.95871,
    19.57063, 20.0078, 20.85755, 21.08295, 20.50464, 19.68516, 19.93076,
    20.95179, 21.63695, 20.37842, 18.72233, 18.89332, 23.52264, 27.02943,
    22.17672, 21.70859, 25.00801, 27.62862, 27.09805, 27.33153, 27.88654,
    27.62548, 21.71112,
  19.013, 18.79254, 19.52046, 20.80572, 21.2957, 20.72658, 20.24549,
    19.96232, 19.7415, 19.94719, 19.75609, 20.90859, 23.02875, 23.40084,
    22.83925, 27.54613, 34.66532, 28.28752, 22.46321, 26.0743, 25.35079,
    20.37998, 21.19549, 22.48596, 25.68583, 26.13164, 25.58623, 38.35979,
    38.94483, 21.58035,
  18.83781, 19.12443, 20.22826, 21.65435, 22.26281, 21.56592, 21.14347,
    22.88902, 23.23903, 23.04043, 23.70617, 23.86412, 23.2544, 22.93994,
    27.58511, 37.01407, 36.55865, 27.0111, 23.68472, 23.95138, 21.90914,
    20.49548, 21.29639, 24.06776, 26.41502, 23.76294, 29.76439, 48.48964,
    42.33219, 19.91838,
  18.96999, 19.42784, 20.67896, 21.95228, 21.77685, 23.24853, 25.84154,
    24.58766, 22.97716, 23.33559, 23.78145, 22.64399, 20.73363, 20.63943,
    24.70085, 29.06367, 26.28123, 23.55371, 22.08714, 21.85005, 21.08787,
    20.65242, 22.13974, 25.35, 25.42261, 22.52729, 36.39016, 49.32995,
    29.64085, 19.8093,
  20.45799, 20.72157, 21.8918, 22.09358, 22.34178, 26.12176, 26.33583,
    22.75538, 22.68292, 23.23227, 22.54463, 20.92676, 19.88582, 23.69442,
    27.37345, 24.02994, 23.34718, 25.42429, 25.25002, 23.05576, 20.58652,
    21.97062, 26.6992, 28.57401, 24.15504, 23.75486, 33.69845, 36.23911,
    22.30694, 19.85573,
  22.7651, 23.39001, 26.05278, 29.31623, 29.1666, 26.45532, 21.9783, 21.2779,
    21.34627, 20.77193, 21.37605, 25.29282, 27.30804, 28.07048, 27.26982,
    26.48733, 27.24109, 28.22824, 27.51122, 25.44333, 24.90054, 26.32462,
    28.6367, 27.29138, 30.1341, 41.17894, 38.21521, 25.12364, 20.75524,
    18.91273,
  29.47715, 36.80631, 37.12934, 29.55558, 29.53155, 29.05796, 25.80632,
    26.83139, 28.04219, 32.28798, 37.97122, 29.53077, 26.55364, 25.71771,
    24.63265, 26.13825, 28.28792, 28.32035, 26.77466, 25.71393, 28.7175,
    29.23496, 26.02047, 23.09802, 28.34483, 36.21611, 30.4988, 20.55914,
    19.33528, 18.50898,
  47.58406, 40.56973, 36.45027, 33.29512, 34.0227, 28.47294, 32.77684,
    33.9792, 29.63573, 34.72933, 36.51258, 23.45823, 24.20523, 25.83483,
    24.96788, 26.02881, 25.63867, 25.44743, 24.61609, 25.15498, 29.09895,
    28.20977, 22.71829, 25.53672, 30.18658, 24.90619, 20.05078, 19.48029,
    19.39741, 18.76156,
  63.20534, 49.03083, 50.0503, 56.25647, 58.20017, 54.69232, 49.97813,
    43.4077, 49.86332, 36.66454, 27.60528, 22.57087, 28.0156, 29.34618,
    27.20091, 25.86422, 26.02728, 25.00914, 23.8698, 27.21782, 30.55505,
    25.88111, 22.20794, 28.86656, 33.57136, 22.50181, 19.22692, 19.68823,
    20.03717, 19.2721,
  71.65591, 60.39828, 61.52653, 66.87576, 69.89372, 70.79314, 63.54527,
    62.83711, 53.84041, 36.21877, 39.27089, 40.01023, 45.75426, 46.99083,
    41.04122, 32.16887, 26.56703, 28.52295, 30.74347, 33.21872, 30.22356,
    26.58877, 30.49356, 28.79752, 25.31847, 20.35311, 19.34386, 19.32194,
    19.9059, 19.39234,
  55.09585, 64.27959, 71.44114, 78.22139, 79.19848, 70.87564, 68.97063,
    72.07533, 49.61855, 48.19094, 56.64021, 54.66698, 48.56058, 43.31915,
    45.73423, 32.56239, 31.24313, 31.83271, 34.43433, 36.06023, 31.23179,
    29.41722, 28.55948, 24.18246, 19.95123, 20.1292, 19.53175, 19.19559,
    19.25211, 18.96392,
  40.56062, 50.65955, 57.2122, 56.87787, 49.801, 50.33153, 57.33196, 43.5374,
    42.70656, 51.28608, 46.00803, 40.01135, 35.17274, 35.17941, 34.95883,
    31.08578, 33.81437, 31.53356, 30.81248, 31.8845, 27.42808, 25.18528,
    22.16509, 20.92731, 20.52302, 20.12788, 19.66653, 19.36755, 19.11864,
    18.75846,
  32.75383, 34.51941, 35.10103, 31.74762, 28.60152, 32.70117, 36.46859,
    31.06906, 35.5163, 39.05592, 30.58707, 28.39321, 32.55734, 30.91203,
    31.05387, 31.42301, 32.31004, 29.30033, 29.06453, 30.48413, 22.99491,
    22.0895, 21.21587, 20.92286, 20.45118, 20.15294, 19.65221, 19.12904,
    19.00005, 18.75336,
  26.89736, 27.01417, 25.07558, 23.90464, 24.40483, 26.15735, 27.16603,
    28.42857, 28.7947, 26.59022, 25.20522, 30.06206, 33.50197, 31.87048,
    37.04955, 35.30254, 30.28386, 26.01741, 29.07763, 29.60669, 21.79337,
    21.75804, 21.32643, 21.03354, 19.98612, 19.82358, 19.57485, 18.84661,
    18.76131, 18.63775,
  25.85792, 25.40302, 22.70804, 21.88666, 22.51649, 23.15339, 24.05121,
    24.37246, 23.45722, 21.899, 25.42515, 29.60621, 27.44409, 29.5456,
    33.78962, 31.90462, 29.93389, 28.1211, 31.54481, 30.13427, 24.0561,
    22.4957, 21.43529, 21.0591, 19.75105, 19.40267, 19.36345, 18.82862,
    18.66443, 18.56063,
  25.74899, 24.7592, 22.3673, 20.75223, 21.20165, 21.46688, 21.73246,
    21.75379, 21.05295, 23.39367, 27.51245, 25.87038, 23.95336, 25.98148,
    27.26781, 26.8829, 28.11384, 29.92343, 30.98409, 30.77174, 27.91786,
    24.93161, 21.7045, 21.12856, 20.09055, 19.41528, 19.23184, 18.8968,
    18.6723, 18.57345,
  24.50541, 23.92775, 21.97305, 20.41724, 20.45735, 20.71637, 20.69581,
    20.39376, 21.10717, 25.3223, 26.72889, 22.68901, 24.02857, 25.23093,
    24.92157, 24.45929, 25.14153, 26.22526, 26.57004, 27.1951, 27.99425,
    27.44749, 23.38626, 21.86965, 20.64468, 19.84139, 19.25812, 18.87299,
    18.67216, 18.57273,
  25.01906, 23.24115, 21.69931, 20.72338, 20.70737, 20.15221, 20.19361,
    20.33111, 22.73667, 26.114, 24.29108, 21.20329, 23.27279, 24.1366,
    23.91368, 23.53918, 23.35386, 23.20927, 23.8027, 24.09159, 25.64224,
    26.52234, 23.86259, 24.22697, 22.58922, 20.53087, 19.34114, 18.95306,
    18.68041, 18.57209,
  25.16261, 23.36583, 21.57593, 20.57859, 21.30193, 21.5492, 21.64578,
    21.38203, 23.83827, 25.42656, 21.9725, 20.78971, 22.1757, 22.8641,
    22.8222, 23.27633, 23.31052, 22.49592, 22.34872, 22.27285, 23.75401,
    24.2233, 22.02993, 24.3347, 24.5657, 21.67444, 19.55538, 19.47505,
    19.03302, 18.61797,
  24.98258, 23.4503, 22.41164, 22.10506, 22.76363, 23.10499, 24.65821,
    26.19855, 27.61306, 24.91153, 20.78834, 21.24916, 22.35407, 23.34346,
    23.46631, 23.82829, 24.23703, 23.28658, 21.98621, 21.9941, 22.87598,
    22.47178, 21.19924, 22.20333, 23.61045, 23.28518, 21.26565, 20.00267,
    19.53533, 18.81504,
  24.7766, 24.72625, 22.75061, 22.2373, 23.59943, 24.99046, 26.10797,
    27.13276, 28.65226, 25.56278, 20.67365, 21.71027, 22.83295, 23.94378,
    24.44274, 24.84989, 24.60179, 23.85937, 22.54519, 21.94789, 22.0777,
    21.76038, 21.66634, 21.30339, 21.17258, 22.77407, 22.72615, 20.94802,
    20.57199, 19.52412,
  25.34484, 26.72687, 25.27135, 24.15662, 24.62077, 25.6116, 27.1195,
    28.56974, 27.27909, 24.46734, 21.1468, 22.18307, 23.59014, 24.25908,
    24.18205, 24.55662, 24.00368, 23.34245, 22.86263, 21.93934, 21.97879,
    22.26689, 21.48302, 20.48145, 20.20632, 21.27178, 22.90446, 22.06869,
    20.74942, 19.62592,
  26.65462, 28.04598, 26.82187, 25.12881, 24.73957, 24.66661, 28.01825,
    29.90368, 25.29705, 22.09682, 21.65776, 22.7627, 23.88408, 24.11996,
    23.85828, 23.74035, 23.26677, 22.97579, 22.6565, 21.73256, 22.03208,
    23.23092, 23.06084, 21.91194, 21.72197, 22.1683, 24.5376, 24.46468,
    20.72398, 18.84028,
  28.92995, 30.71816, 25.55672, 24.42718, 25.1521, 25.42157, 27.73468,
    27.44007, 22.3873, 20.93649, 21.66626, 22.704, 23.33332, 23.61938,
    24.17894, 23.98668, 23.00771, 22.5424, 22.73792, 23.04861, 23.82373,
    24.46162, 23.89811, 22.98557, 22.88171, 23.25967, 24.43199, 26.49054,
    24.09058, 19.56114,
  27.58301, 25.9498, 24.87258, 28.36368, 28.85352, 28.23504, 28.34, 24.57466,
    21.03393, 21.02419, 20.93912, 21.14248, 21.65107, 22.42252, 23.74522,
    24.23447, 23.89846, 23.93719, 23.7627, 23.51991, 23.89544, 23.48373,
    22.1617, 21.45764, 21.88755, 22.66184, 23.03551, 23.78513, 24.12941,
    20.78507,
  25.98221, 24.89547, 26.694, 29.56036, 29.13884, 29.69589, 29.38964,
    24.29139, 20.76751, 21.32286, 21.51796, 22.18328, 23.05202, 23.71804,
    24.56723, 25.16828, 24.64633, 23.63799, 22.93681, 21.95856, 21.37589,
    21.14841, 20.71507, 20.49575, 20.79036, 21.58751, 22.00077, 21.26402,
    20.70337, 19.40896,
  18.4803, 18.55455, 18.62431, 18.66916, 18.65058, 18.64763, 18.66314,
    18.7097, 18.74777, 19.03045, 20.59759, 21.05286, 18.99147, 19.32765,
    19.62516, 18.93233, 18.76858, 18.80552, 18.84178, 19.59631, 20.26245,
    19.75422, 19.87062, 20.75937, 21.68793, 22.2647, 26.6943, 30.66924,
    24.08369, 20.83715,
  19.02847, 19.22309, 18.87092, 19.37426, 19.08106, 18.75369, 18.84349,
    18.92911, 19.13346, 19.62096, 20.66382, 21.62856, 21.88722, 20.88772,
    20.04667, 20.203, 19.16556, 19.33301, 20.39896, 21.49204, 21.1892,
    20.14087, 20.2802, 23.30945, 30.33822, 34.28041, 32.09206, 38.82688,
    26.66168, 22.3762,
  19.07343, 19.14924, 19.04549, 19.13348, 18.90169, 18.74191, 18.79583,
    18.99783, 19.25137, 19.47771, 19.78802, 20.61482, 21.38074, 21.93996,
    21.97812, 20.35851, 20.21705, 21.24771, 21.30194, 21.6307, 23.16124,
    25.3647, 27.11132, 30.31804, 38.95632, 46.30587, 38.52535, 38.03296,
    26.12141, 23.51609,
  19.00223, 19.04621, 19.33282, 19.61525, 20.01355, 20.8928, 20.9135,
    20.29867, 20.34546, 20.85171, 21.305, 21.82874, 21.58361, 21.09201,
    22.98978, 24.77594, 23.96797, 21.44327, 21.13707, 22.36691, 28.34018,
    32.72117, 30.62082, 38.65962, 45.68192, 40.86321, 45.15868, 35.06942,
    25.46844, 21.50322,
  19.89903, 19.17594, 19.70304, 20.33076, 21.20719, 21.6363, 21.28511,
    20.9617, 22.12683, 23.37577, 22.93263, 22.07357, 21.34365, 22.03277,
    23.5961, 24.23416, 22.36786, 20.53165, 22.93058, 31.47204, 37.14967,
    29.55495, 29.73909, 34.0744, 36.2413, 35.29873, 34.52237, 36.92681,
    34.91623, 24.53724,
  19.68358, 19.821, 21.45813, 24.07091, 24.3196, 22.59828, 22.3481, 21.65794,
    21.29341, 21.41047, 21.40209, 24.18254, 28.8155, 30.05432, 33.20416,
    39.51035, 44.80107, 38.71593, 31.57388, 35.9217, 33.11869, 25.68959,
    27.69287, 30.28712, 34.44079, 34.94865, 35.38264, 54.95275, 51.30954,
    24.39697,
  19.87885, 21.16474, 23.40762, 25.55488, 25.28413, 24.09263, 25.50715,
    28.94234, 29.28644, 28.62724, 30.45679, 30.58898, 29.32521, 30.98776,
    38.73878, 48.83166, 46.49297, 37.44419, 31.26724, 31.04338, 27.41078,
    25.11686, 27.17205, 32.53045, 36.98093, 36.4558, 44.89492, 61.92366,
    51.02688, 21.07318,
  20.56166, 22.28764, 24.59427, 26.46646, 26.39282, 30.40082, 35.98741,
    32.5881, 28.93549, 29.24505, 29.19385, 27.55035, 25.65629, 27.98907,
    33.49313, 37.53448, 34.80412, 31.67477, 27.01343, 26.45679, 25.00218,
    24.68926, 28.26238, 34.14177, 35.41351, 34.72199, 49.53229, 61.47854,
    38.06969, 20.64215,
  22.95062, 23.57125, 26.5068, 27.95126, 28.90145, 34.1398, 33.22263,
    28.87714, 29.26982, 28.83446, 27.06468, 24.98159, 25.41516, 33.8284,
    40.56238, 33.19436, 30.59913, 32.94705, 32.70227, 28.77137, 25.0343,
    28.83333, 37.28735, 40.33164, 32.89022, 34.61978, 47.16703, 49.00458,
    27.33562, 20.62587,
  28.77766, 35.20551, 37.32401, 38.47791, 38.63847, 34.88118, 25.49008,
    25.1147, 24.60422, 24.62426, 28.21821, 37.09264, 40.97476, 40.21308,
    36.25101, 34.87771, 36.26615, 37.47839, 34.92128, 30.5951, 31.13779,
    33.68464, 36.71515, 37.5941, 45.2842, 58.75872, 51.8492, 29.76694,
    21.57932, 19.10969,
  42.18568, 49.11091, 48.63061, 42.42083, 42.82943, 38.62399, 30.57573,
    34.07556, 38.62351, 46.40748, 54.41138, 40.70431, 35.27445, 33.08372,
    31.03021, 33.19923, 35.90504, 35.11, 32.38536, 30.67993, 34.36865,
    35.3866, 31.28801, 29.43538, 36.80899, 43.87447, 34.2985, 20.47431,
    19.63087, 18.58425,
  61.56117, 50.0891, 48.07553, 48.12213, 47.12189, 38.91289, 46.00187,
    49.60323, 46.57975, 49.36999, 46.31206, 31.35656, 31.97679, 33.45211,
    32.53647, 33.91971, 32.83304, 31.49537, 29.92481, 31.26156, 34.93787,
    33.06626, 26.1554, 30.8051, 37.13743, 28.30078, 20.71073, 19.94654,
    19.83974, 18.94699,
  75.36532, 62.85073, 72.19099, 80.05682, 81.15349, 75.80109, 66.56094,
    52.24825, 53.2067, 43.35984, 34.85233, 29.0378, 36.78082, 41.75692,
    38.5591, 34.44705, 33.53523, 31.07138, 29.48232, 36.6015, 39.68998,
    29.4652, 26.40443, 34.08925, 38.07454, 23.76594, 19.46951, 20.34495,
    20.65348, 19.61624,
  83.07967, 94.07847, 96.3987, 98.32548, 91.96355, 86.65847, 80.02772,
    73.19741, 57.74089, 46.51683, 55.67363, 57.84466, 63.87189, 64.87256,
    56.96179, 43.43034, 34.30099, 36.33856, 39.71242, 43.05784, 37.31877,
    30.24328, 36.97769, 32.33475, 25.87697, 20.95131, 19.82973, 19.7648,
    20.38177, 19.72469,
  79.77749, 79.68049, 82.40392, 79.95354, 71.72462, 71.70734, 84.45808,
    79.94418, 66.0713, 70.11834, 74.25679, 65.63821, 59.57743, 64.28989,
    62.05708, 45.30147, 42.43353, 44.46529, 49.4282, 49.82608, 39.71183,
    37.6188, 34.10503, 25.19941, 20.40867, 20.72735, 19.96592, 19.50778,
    19.51033, 19.12914,
  73.75085, 73.7141, 72.31062, 67.17565, 68.30066, 74.57956, 82.76272,
    88.66384, 70.74429, 62.93553, 62.83154, 53.38098, 47.70166, 54.398,
    50.5836, 45.89974, 47.82185, 45.21711, 46.15785, 45.94907, 34.09565,
    29.6519, 24.8737, 21.97486, 21.26945, 20.72464, 20.01715, 19.67148,
    19.31868, 18.885,
  65.29132, 61.17634, 55.69811, 53.81673, 55.64144, 55.75958, 60.97506,
    68.92603, 54.324, 51.12418, 46.35141, 44.41973, 50.64882, 49.7509,
    46.985, 46.73997, 45.84644, 40.57923, 41.34543, 41.74934, 26.09648,
    23.22153, 22.42148, 22.42365, 21.29844, 20.70195, 20.05014, 19.36322,
    19.16581, 18.90203,
  50.13593, 46.59776, 42.17871, 42.30154, 43.37931, 46.69802, 50.13966,
    49.15854, 44.44292, 41.20477, 41.07419, 49.40472, 53.24737, 53.18042,
    55.9216, 50.88467, 41.79404, 36.33642, 41.11315, 38.04407, 23.38329,
    23.83054, 23.39392, 22.66192, 20.57074, 20.31064, 19.98636, 18.97964,
    18.88523, 18.74909,
  43.91831, 42.38968, 36.89301, 35.41712, 38.88343, 42.7944, 42.37531,
    39.12139, 35.80802, 34.37218, 41.86947, 49.65823, 46.38596, 49.46799,
    50.48877, 43.30684, 40.45532, 42.44798, 45.89487, 39.22477, 27.88962,
    26.44292, 24.33372, 22.6019, 20.17878, 19.8339, 19.68192, 18.95306,
    18.76659, 18.6622,
  41.46754, 40.54866, 34.66146, 32.58894, 36.20958, 37.30433, 34.60752,
    31.87394, 30.84282, 38.16132, 47.16204, 44.71642, 42.59597, 43.59586,
    40.41446, 35.73996, 36.73982, 42.45593, 44.60188, 42.19922, 36.20479,
    30.36388, 24.69178, 22.70892, 20.76224, 19.93651, 19.59131, 19.0891,
    18.76555, 18.67422,
  38.7673, 37.99001, 33.0359, 31.53707, 33.2085, 32.46495, 29.84446,
    28.90761, 32.6922, 43.10604, 46.18104, 39.13443, 40.82942, 38.94609,
    34.88468, 32.60323, 33.85994, 37.1316, 39.04636, 39.29526, 36.62113,
    32.76158, 27.19257, 23.76475, 21.53747, 20.56976, 19.65839, 19.11063,
    18.80077, 18.68198,
  38.8195, 36.35057, 32.24803, 31.4584, 31.19767, 28.7272, 28.20703,
    29.82719, 36.92491, 44.01155, 40.09431, 35.06182, 36.7987, 34.04749,
    31.67616, 31.42845, 32.71686, 33.88845, 34.80145, 34.208, 32.82035,
    31.43969, 28.67539, 27.8957, 24.88061, 21.66348, 19.7905, 19.24814,
    18.83595, 18.69604,
  37.75896, 36.29848, 31.41604, 29.70078, 30.32089, 30.38152, 31.21424,
    32.61279, 38.71092, 41.5858, 34.1996, 31.77141, 31.99404, 30.54708,
    29.6278, 31.12484, 32.92058, 32.21675, 31.20519, 29.79421, 29.59318,
    29.22783, 26.99994, 28.96564, 28.42304, 23.52615, 20.18989, 20.07983,
    19.32534, 18.75097,
  37.22155, 35.459, 32.98001, 31.97193, 32.63183, 33.92512, 36.67786,
    37.50828, 41.77726, 39.74352, 30.93165, 30.59727, 30.81323, 31.10428,
    31.6007, 33.33868, 34.5345, 32.51217, 29.52455, 27.99916, 27.52316,
    26.88639, 25.90716, 26.86834, 27.8657, 26.26066, 22.8588, 20.81177,
    19.97066, 19.01564,
  35.88628, 37.71933, 32.91544, 31.94817, 33.80128, 35.17636, 37.01441,
    38.23808, 43.04486, 39.36046, 29.47802, 30.53992, 31.58352, 33.31089,
    34.87493, 36.15179, 34.98739, 32.37205, 28.67311, 25.92762, 26.13955,
    26.56396, 25.95129, 24.56433, 23.76451, 25.3175, 24.84411, 22.05974,
    21.30719, 19.97074,
  37.87394, 41.29963, 36.69068, 34.51905, 35.12379, 35.67091, 37.38816,
    40.27972, 41.97401, 36.16393, 29.80961, 31.54387, 33.98735, 35.62776,
    35.79599, 35.68084, 33.37238, 30.47779, 27.22927, 24.59064, 26.25571,
    27.39519, 24.80959, 22.08064, 21.40414, 23.03229, 25.018, 23.67897,
    21.6563, 20.20084,
  41.21577, 44.03945, 39.3336, 35.91153, 36.43589, 35.42624, 38.30606,
    41.00488, 38.74066, 31.85419, 30.97141, 33.54974, 35.94403, 36.35507,
    35.2366, 33.6834, 31.11095, 28.57506, 26.01163, 24.11134, 26.13755,
    28.20389, 26.46233, 23.87406, 23.39306, 24.32616, 27.34782, 27.03367,
    21.74133, 19.15004,
  44.18539, 45.66745, 38.17004, 36.29811, 38.98529, 38.53343, 40.69434,
    39.95511, 33.58709, 30.31116, 32.09828, 34.88802, 36.26376, 35.79292,
    34.96354, 32.88004, 29.48021, 27.03311, 25.83213, 25.94326, 28.80942,
    30.30358, 27.84489, 25.59904, 25.01304, 25.88035, 27.50383, 29.74128,
    26.22454, 20.11605,
  40.13984, 35.87741, 34.51314, 39.40114, 41.87149, 44.17922, 43.49878,
    36.76054, 30.51814, 31.05472, 32.03632, 33.15217, 33.58929, 33.51984,
    33.66736, 32.30298, 30.09434, 29.04489, 27.55242, 26.87166, 28.60541,
    27.96198, 25.00748, 23.40795, 23.79614, 24.98705, 25.55365, 26.36462,
    26.38093, 21.90096,
  35.91904, 34.41341, 37.23439, 39.68576, 39.4063, 43.29106, 44.99344,
    36.02828, 30.36063, 32.45614, 33.62852, 34.90842, 35.38925, 34.99841,
    34.53929, 33.83917, 31.21544, 28.45721, 26.32692, 24.51953, 23.91834,
    23.06985, 22.13069, 21.78476, 22.29662, 23.34215, 23.80965, 22.83622,
    21.86072, 19.95515,
  24.83862, 25.02131, 25.32184, 25.6199, 25.66899, 25.82798, 26.12306,
    26.58948, 27.19651, 28.42776, 30.86528, 31.01825, 26.83797, 27.68079,
    27.92679, 26.64323, 26.70305, 27.50992, 28.78004, 31.24185, 32.82319,
    31.66665, 33.01596, 36.58401, 40.29159, 43.2187, 51.27982, 55.13126,
    34.87735, 28.51601,
  26.5147, 27.131, 26.4087, 27.67526, 27.06713, 26.6337, 27.2611, 27.83647,
    28.60763, 29.65449, 31.2135, 32.99746, 33.76366, 31.27129, 29.47101,
    30.35223, 29.04476, 31.11418, 34.25718, 37.08413, 37.93728, 39.24181,
    43.16676, 51.76311, 60.6666, 59.48625, 54.51974, 58.50692, 36.54892,
    30.60097,
  24.28245, 24.43822, 24.66459, 24.98914, 25.04064, 25.35354, 25.63169,
    26.17454, 26.92344, 27.76947, 28.9284, 30.7896, 32.48776, 34.30538,
    35.47916, 33.80524, 36.26675, 40.50703, 43.77778, 49.60765, 58.4099,
    67.97976, 73.11266, 75.66351, 77.15077, 72.28094, 65.28379, 54.60042,
    36.88967, 32.60365,
  24.07177, 24.84134, 26.50665, 28.42084, 30.19962, 32.22305, 32.21423,
    31.30959, 32.32783, 34.02591, 35.03532, 35.99265, 36.81934, 37.8936,
    44.15443, 49.26608, 48.97884, 48.09903, 54.9108, 63.15157, 75.68222,
    81.35904, 75.86958, 82.04202, 81.97963, 78.41946, 70.96387, 51.64108,
    36.07442, 29.29628,
  27.71841, 27.04535, 29.87838, 31.97478, 33.71551, 33.54334, 32.80978,
    32.87626, 34.83218, 36.20821, 35.35143, 36.22688, 38.22891, 42.95848,
    48.27088, 52.8454, 54.03587, 54.12962, 61.00484, 72.07123, 76.31729,
    64.23779, 64.66109, 71.80392, 77.36013, 76.16327, 66.80881, 70.12699,
    61.55569, 36.98707,
  28.77737, 31.23488, 35.16121, 39.02652, 37.61214, 33.78323, 33.86303,
    33.9419, 34.94283, 39.04827, 46.00011, 58.25076, 71.96111, 74.32895,
    78.98089, 85.66037, 91.2131, 84.09451, 73.39433, 72.97321, 64.75517,
    56.03624, 62.62416, 69.87177, 77.85333, 77.24718, 71.44298, 84.77898,
    75.2481, 35.97434,
  30.95965, 34.85319, 39.71553, 44.89339, 47.20329, 50.5378, 59.11023,
    69.4047, 73.4749, 75.375, 78.59167, 76.24524, 69.80579, 72.40783,
    75.8784, 79.08199, 78.35472, 71.46877, 60.94799, 61.61583, 58.33972,
    58.967, 66.30805, 75.65477, 77.73314, 68.23251, 70.00076, 80.07389,
    65.06509, 28.56082,
  36.34303, 43.21524, 51.25207, 59.90791, 65.42541, 76.14555, 84.04873,
    70.86384, 61.73781, 62.37036, 58.75587, 53.96201, 49.52686, 50.93206,
    53.49681, 57.88599, 59.86038, 58.06866, 51.71886, 54.15589, 54.86154,
    58.86504, 67.56776, 74.41693, 70.25788, 64.98369, 76.02965, 76.69349,
    52.70346, 28.88891,
  50.23222, 56.38755, 63.18892, 67.22731, 68.35676, 71.43197, 61.65298,
    54.65755, 55.54589, 54.40355, 52.2017, 51.70234, 55.90368, 69.48871,
    77.2348, 60.91383, 62.13203, 68.23712, 68.36874, 62.59827, 60.71072,
    74.70941, 89.57417, 89.4823, 74.13941, 80.90137, 84.4099, 69.5631,
    37.81371, 28.53106,
  73.29972, 83.06104, 80.26629, 82.63736, 73.88229, 60.86506, 43.34944,
    50.52136, 53.9605, 63.56995, 76.33544, 90.45489, 89.19147, 84.41689,
    76.17501, 80.72772, 86.20596, 86.33542, 82.11696, 80.59324, 90.0379,
    93.25967, 90.86785, 80.70714, 87.84689, 101.1231, 83.3248, 47.63403,
    28.6818, 25.25355,
  96.72122, 91.74387, 87.22882, 75.25692, 83.78717, 84.30444, 82.63681,
    92.74329, 102.4924, 107.915, 99.84001, 73.72343, 67.84792, 66.40461,
    68.50539, 75.5995, 81.67039, 82.28218, 80.7291, 83.06422, 95.29432,
    92.67063, 73.06953, 64.81422, 72.79208, 72.4287, 49.16255, 28.80632,
    27.00423, 24.82828,
  97.88849, 78.5612, 87.78448, 97.17247, 100.9606, 92.50809, 98.93246,
    95.99309, 85.8835, 73.50147, 62.26329, 54.46321, 60.30326, 66.36521,
    69.81725, 72.27089, 72.34122, 72.51384, 70.88875, 73.77264, 83.74168,
    77.65008, 59.30887, 67.77596, 70.83957, 49.46814, 28.1596, 29.21885,
    27.99066, 25.85763,
  112.9938, 113.3995, 118.286, 120.7226, 121.521, 118.3855, 99.34308,
    83.66977, 83.51624, 59.9637, 57.76448, 60.90368, 73.15041, 82.32054,
    80.28779, 69.66239, 70.86007, 68.29725, 66.90807, 74.72124, 79.58743,
    68.94666, 61.12726, 60.00178, 54.44189, 38.16545, 28.53398, 31.07791,
    30.07156, 27.58718,
  118.7323, 121.2763, 121.6343, 119.6927, 116.4485, 112.9848, 110.7074,
    110.5285, 91.68207, 92.65205, 108.2659, 103.2868, 110.7083, 113.9342,
    97.47952, 80.68672, 80.62192, 87.0816, 93.93964, 92.23341, 79.57578,
    64.81587, 59.08215, 45.2998, 36.44548, 32.77346, 29.82251, 29.00704,
    28.88425, 27.44884,
  116.3893, 112.9411, 106.8043, 101.6191, 99.63386, 104.9176, 113.2027,
    114.5087, 111.5997, 112.7283, 112.5172, 108.9595, 112.5536, 112.6383,
    108.1089, 107.9546, 100.8651, 101.8635, 103.1209, 92.40903, 62.91882,
    55.25204, 42.81879, 35.55089, 32.74998, 31.64642, 29.30891, 27.68686,
    26.73298, 25.88883,
  102.9116, 99.44765, 99.56639, 100.4347, 104.0412, 112.8086, 115.7758,
    114.2286, 110.3899, 108.0642, 106.4136, 98.69785, 95.87675, 109.7914,
    107.9119, 105.2853, 103.3921, 90.91549, 81.76576, 68.18899, 45.1319,
    42.35813, 35.00592, 33.61959, 32.71944, 30.68782, 28.47235, 27.43254,
    26.2919, 25.50314,
  89.21758, 83.69075, 86.44725, 91.22477, 96.50709, 101.2234, 104.1413,
    104.0984, 100.3699, 96.50745, 87.86501, 98.50725, 114.2171, 110.0344,
    103.7313, 96.44981, 85.76682, 72.64151, 67.14082, 60.56168, 38.43675,
    39.37908, 35.34951, 33.64645, 31.74439, 30.52789, 28.22058, 26.39847,
    25.80963, 25.46819,
  71.6893, 74.33122, 76.23485, 80.81789, 84.10033, 87.19917, 88.47163,
    89.42421, 89.31686, 88.08301, 101.3265, 115.7558, 115.9645, 115.2746,
    113.8214, 91.48505, 67.73656, 58.83615, 64.02945, 58.14114, 38.92575,
    39.99073, 36.33163, 34.19174, 30.66908, 29.25528, 27.88347, 25.55076,
    25.31072, 25.07006,
  78.25032, 78.29696, 70.94797, 68.52382, 70.58518, 71.46632, 73.58648,
    77.45761, 81.25754, 91.86359, 110.9115, 114.3671, 96.19643, 94.69742,
    85.39749, 73.69247, 72.19358, 76.68314, 79.03829, 67.10329, 47.47509,
    41.96944, 36.95065, 33.9576, 29.5472, 27.87921, 26.95911, 25.49446,
    25.13435, 24.9871,
  79.39314, 74.32691, 63.85246, 57.22807, 59.03912, 61.17358, 66.01288,
    73.08397, 83.31696, 99.41815, 105.1202, 83.74907, 74.10474, 70.77557,
    64.35098, 62.96634, 69.33604, 77.86256, 78.12085, 71.30534, 58.20601,
    46.47767, 37.73542, 34.40172, 30.8552, 28.08989, 26.93637, 25.75802,
    25.12385, 25.03817,
  71.49595, 64.72937, 54.44047, 49.84059, 52.80368, 57.95878, 64.59829,
    72.42822, 81.62857, 89.33885, 80.07265, 61.1705, 65.07682, 63.6738,
    60.99356, 60.90574, 64.51406, 66.57495, 65.85546, 61.63408, 55.61721,
    51.67994, 43.8187, 37.73906, 33.38309, 29.80002, 27.03603, 25.81451,
    25.16376, 25.07888,
  67.93315, 57.09918, 50.95037, 49.48047, 53.87105, 57.06202, 64.25187,
    69.10809, 75.76062, 76.29082, 61.67353, 52.94054, 59.07646, 59.49737,
    59.03109, 58.9857, 57.74879, 55.51366, 54.021, 51.75948, 50.25481,
    48.82799, 47.03797, 45.40888, 38.9509, 31.12948, 27.09566, 26.10112,
    25.20862, 25.0527,
  62.77833, 55.74925, 49.18259, 49.64181, 58.75658, 64.39516, 66.95943,
    65.22245, 66.55141, 62.7121, 48.72672, 49.76305, 54.12241, 56.0117,
    55.16331, 55.05808, 52.68074, 47.74365, 45.77957, 45.43341, 45.58142,
    45.07017, 43.28338, 44.35834, 43.23621, 34.49475, 28.62322, 28.29749,
    26.52751, 25.17692,
  63.68399, 59.70379, 59.49202, 64.08496, 70.21616, 71.08394, 72.93918,
    69.61449, 69.00838, 58.69685, 46.4285, 52.89603, 56.76597, 59.51817,
    57.81757, 55.30134, 52.42188, 47.83614, 44.23912, 43.88454, 43.58169,
    42.20166, 40.7603, 40.62424, 41.37126, 39.77643, 34.37085, 29.72782,
    27.97704, 25.91629,
  65.36047, 67.26796, 64.2388, 67.38652, 71.63721, 70.35185, 67.38099,
    65.93044, 69.47431, 60.13915, 47.42261, 55.31071, 59.05985, 61.46745,
    59.34738, 56.6812, 52.38572, 48.78938, 45.49636, 42.71292, 42.71446,
    42.59766, 40.2453, 37.79236, 37.07098, 39.56562, 39.33556, 33.89357,
    31.30744, 28.48625,
  75.14896, 80.9271, 79.44533, 75.28981, 71.73021, 67.87108, 69.85201,
    73.34422, 69.09314, 57.04258, 53.55708, 59.99252, 63.03212, 61.43507,
    56.12696, 53.61358, 50.90114, 48.59555, 46.58215, 43.56434, 43.42062,
    42.36908, 38.17539, 35.33421, 35.89768, 38.5264, 41.24041, 38.1066,
    31.65637, 28.53369,
  86.53972, 90.47035, 81.13062, 73.22151, 68.8094, 65.18427, 71.6103,
    72.44022, 61.33459, 53.53118, 58.50724, 61.82723, 61.50607, 57.67028,
    53.72717, 51.78365, 49.62537, 47.51229, 45.16533, 42.34044, 43.39817,
    45.88538, 45.14701, 42.4548, 42.74186, 44.88115, 48.48647, 45.25346,
    32.3107, 26.18707,
  91.98058, 87.52931, 77.29565, 74.35698, 74.30783, 72.70464, 74.80122,
    67.73921, 54.65675, 56.49414, 60.46271, 60.77042, 58.88555, 55.75407,
    54.73598, 51.90091, 47.40484, 45.65411, 47.14502, 49.44357, 51.9417,
    52.53587, 48.93198, 46.96012, 47.29932, 49.30841, 50.43929, 51.65785,
    43.87175, 29.44289,
  79.18803, 73.58018, 76.33305, 82.96425, 84.2254, 85.12329, 76.76781,
    60.90337, 52.97224, 55.47636, 52.61466, 50.31957, 49.6778, 50.29116,
    52.28098, 52.51573, 52.14807, 53.69519, 53.45956, 52.1469, 52.0646,
    49.59858, 45.60574, 44.15221, 45.42033, 46.89294, 46.50499, 44.16505,
    41.01129, 33.1258,
  75.30959, 77.96376, 80.76225, 80.67865, 80.65238, 85.79042, 82.37061,
    62.76625, 52.98173, 55.97021, 56.40875, 58.9454, 60.96665, 61.25956,
    60.60924, 59.66567, 55.61463, 50.88997, 48.77812, 46.25431, 43.72551,
    42.14969, 40.79732, 40.24059, 40.39796, 40.67713, 39.42574, 35.16344,
    31.19431, 26.67309,
  31.24426, 31.4346, 31.73112, 32.04766, 32.23407, 32.55486, 32.97291,
    33.55786, 34.32583, 35.6353, 37.85943, 38.34444, 35.94627, 37.59668,
    38.68594, 38.62191, 39.63807, 41.09892, 42.67658, 45.06314, 46.42303,
    45.52574, 46.61449, 49.48902, 51.72254, 52.33934, 56.82441, 57.63,
    41.22523, 35.45488,
  31.89548, 32.18395, 31.62265, 32.62968, 32.3378, 32.36649, 33.33819,
    34.38794, 35.78749, 37.57286, 39.98825, 42.95377, 45.18293, 44.66258,
    44.68512, 46.1153, 45.5675, 47.18748, 49.26248, 51.15187, 51.70504,
    52.17657, 53.7303, 58.1058, 62.37333, 58.46676, 52.25712, 55.92005,
    41.78101, 37.05367,
  29.64494, 30.04926, 30.76352, 31.57018, 32.52027, 33.83876, 35.36656,
    37.44634, 39.90835, 42.58488, 45.68783, 49.33185, 52.76995, 56.05995,
    57.92831, 56.94336, 58.46369, 60.79801, 62.80857, 66.87705, 73.16573,
    78.74603, 78.97354, 76.10353, 73.35709, 68.80605, 61.66279, 52.94198,
    41.38082, 38.12822,
  33.84009, 35.51166, 37.95565, 40.59023, 43.07685, 45.82362, 47.36235,
    48.59977, 51.31152, 54.29853, 56.65689, 58.71253, 59.81816, 60.34448,
    64.2835, 66.6119, 64.27126, 62.34432, 66.9659, 72.48173, 80.67961,
    81.49176, 75.69368, 79.43197, 77.51603, 75.41959, 70.90717, 55.75152,
    42.69784, 36.08414,
  38.11444, 38.70388, 42.12238, 45.07558, 47.58871, 49.08014, 50.7103,
    52.82713, 56.09464, 58.41897, 59.08492, 61.37437, 62.98225, 64.44582,
    66.46917, 68.76965, 67.56339, 65.02203, 69.23642, 76.98545, 77.66396,
    67.70821, 68.8865, 75.13219, 80.47382, 80.73112, 75.87377, 79.91801,
    70.52362, 45.3081,
  43.71, 49.40777, 55.50308, 61.58369, 63.24914, 64.12138, 68.36877,
    70.93789, 72.99935, 76.8825, 82.7379, 93.1654, 102.8684, 101.143,
    102.6058, 104.2814, 100.519, 90.88516, 80.00331, 77.41404, 69.49625,
    61.74099, 67.24798, 72.07721, 77.52483, 77.15482, 75.24521, 87.42146,
    78.25935, 41.63491,
  60.24196, 68.4254, 75.05869, 81.60141, 84.91088, 88.85999, 96.65173,
    103.0013, 101.376, 95.74056, 91.40397, 83.01579, 73.57069, 74.23241,
    74.81528, 75.8652, 74.91617, 69.36568, 62.29863, 63.02342, 60.85613,
    60.48996, 64.67484, 70.11371, 70.58971, 65.4862, 68.93723, 76.58113,
    63.61378, 33.93523,
  67.36578, 72.95837, 77.44454, 81.51792, 82.85928, 87.96589, 88.82046,
    72.05129, 62.80025, 62.00684, 58.61637, 55.97374, 54.43245, 56.30667,
    58.52201, 62.05446, 64.77058, 63.52428, 59.54796, 60.94663, 62.07838,
    65.41219, 70.6669, 73.64319, 70.4428, 69.38422, 76.56541, 74.60302,
    54.7199, 35.35734,
  69.28967, 71.21262, 73.68507, 74.49387, 75.037, 76.86086, 68.09381,
    66.85123, 70.8551, 72.39249, 73.42558, 74.9519, 79.21049, 89.42676,
    93.60725, 82.62372, 82.67661, 85.17458, 83.49893, 77.96164, 76.53571,
    84.67368, 91.90741, 88.21516, 77.15784, 81.10016, 79.64557, 64.94794,
    39.34048, 35.2324,
  85.85503, 93.59331, 87.46292, 88.04663, 88.15553, 82.82878, 69.91386,
    79.79799, 83.54472, 90.78462, 99.0753, 107.907, 106.8795, 104.5642,
    101.6114, 105.8814, 106.0729, 101.4023, 95.37865, 93.57722, 95.15688,
    91.26255, 84.92195, 74.78958, 77.86757, 84.8003, 72.42583, 46.90618,
    34.37664, 32.60526,
  116.2423, 116.5001, 113.1767, 102.2213, 109.745, 105.3072, 99.32462,
    105.3866, 109.2528, 105.8354, 93.88496, 77.4369, 74.90776, 75.12947,
    75.07055, 76.23766, 77.14427, 75.92132, 75.02666, 77.80681, 85.37638,
    79.08132, 64.46048, 60.66827, 66.0143, 63.15918, 46.15582, 34.57275,
    34.82404, 32.70241,
  119.1416, 112.6876, 118.0588, 120.1756, 114.3638, 97.11966, 97.48949,
    91.91937, 83.52133, 74.73942, 69.48425, 66.75523, 69.6745, 70.23347,
    67.27074, 65.3652, 63.29816, 63.22232, 63.78229, 68.45433, 76.70599,
    73.95672, 62.60439, 70.63687, 71.85068, 54.74583, 35.66104, 39.25359,
    35.8651, 33.92513,
  126.5913, 126.6181, 128.6234, 129.8752, 129.3265, 126.1466, 114.1693,
    98.98271, 104.6502, 86.63946, 82.40793, 79.32898, 86.07527, 88.52657,
    80.0005, 67.38618, 68.2508, 67.17492, 67.51752, 73.10016, 75.70473,
    68.46394, 61.38377, 57.19861, 54.98037, 46.83909, 37.9179, 39.41118,
    38.44487, 35.49918,
  121.2595, 121.2484, 121.3422, 121.0115, 120.3788, 120.183, 120.6464,
    121.3222, 120.0649, 120.6139, 122.124, 121.1276, 121.9532, 120.5186,
    105.3945, 86.26893, 82.16498, 84.99989, 86.2285, 79.42876, 68.63285,
    59.08036, 52.93827, 43.97948, 39.36098, 38.49791, 36.32277, 35.57868,
    36.00573, 34.9275,
  107.3758, 104.2886, 109.8419, 113.9042, 117.7983, 119.4342, 121.8279,
    122.327, 121.1441, 121.5798, 114.8925, 106.9018, 106.0974, 106.5339,
    103.5083, 98.81201, 87.11484, 81.46301, 79.02343, 71.4576, 53.53922,
    51.71722, 43.9201, 40.67642, 39.45262, 37.76808, 36.05905, 34.60558,
    33.75459, 33.28608,
  106.0989, 111.5984, 114.4417, 116.228, 116.5683, 119.1998, 122.5253,
    115.588, 103.7147, 96.33399, 92.58356, 85.14098, 80.81214, 87.36103,
    83.62776, 79.56274, 77.87503, 68.61528, 64.94879, 57.75791, 45.06886,
    46.57123, 41.85863, 40.38851, 39.41365, 37.68735, 35.80504, 34.91782,
    33.92796, 33.26449,
  94.57892, 92.36766, 94.01934, 96.73668, 99.37166, 101.7033, 102.4478,
    100.8302, 96.31679, 88.07817, 79.12061, 85.46452, 92.77437, 84.41757,
    77.86977, 73.08406, 67.19405, 62.86312, 63.10175, 58.09597, 45.13181,
    46.76768, 42.81786, 40.35344, 38.93123, 37.91473, 35.37803, 33.61697,
    33.3434, 33.10095,
  80.53471, 84.15038, 85.82761, 90.42043, 93.46642, 95.53237, 95.363,
    94.62159, 92.59505, 89.91727, 96.89011, 103.7173, 98.0898, 93.89252,
    87.85262, 75.0369, 64.84057, 62.77599, 66.46104, 59.9902, 45.41137,
    45.60981, 42.68457, 40.91848, 37.51471, 36.29125, 35.2922, 33.01959,
    32.90892, 32.7664,
  93.25562, 91.04758, 83.83271, 80.34917, 81.21075, 79.11189, 77.23933,
    76.28749, 75.57707, 78.89146, 85.69448, 83.17995, 74.55727, 77.83882,
    78.11053, 80.58007, 86.45235, 91.73328, 88.25862, 75.47563, 56.14566,
    48.11741, 43.52969, 41.00932, 37.34124, 35.68497, 34.81524, 33.38207,
    32.8716, 32.79054,
  93.14736, 87.7524, 76.77767, 68.22054, 66.88714, 64.89433, 64.97365,
    67.23607, 71.75392, 80.40366, 81.8442, 71.18845, 71.16356, 71.3512,
    70.15541, 69.77159, 74.09846, 79.49141, 79.76037, 74.8197, 65.78297,
    55.49712, 47.00266, 43.82644, 40.46995, 36.93664, 35.25904, 33.71009,
    32.88053, 32.82254,
  86.94607, 79.0295, 66.93352, 59.19325, 58.22134, 59.25641, 61.848,
    65.52045, 70.69273, 75.35593, 70.35193, 61.25336, 65.56906, 64.10301,
    60.84825, 58.42315, 59.14835, 60.60354, 62.29108, 63.04476, 63.0961,
    62.3634, 55.39716, 48.43427, 43.50613, 38.35265, 35.02396, 33.74073,
    32.94782, 32.8514,
  83.53041, 72.73503, 62.83163, 57.88536, 58.94626, 58.98164, 62.55364,
    64.80587, 69.01607, 68.12466, 56.78036, 51.58811, 53.71015, 53.16603,
    51.40405, 50.87444, 50.41238, 51.17676, 53.38151, 54.85213, 55.82535,
    56.00463, 56.66445, 55.2218, 48.24534, 39.51758, 35.61636, 34.53641,
    33.21972, 32.82032,
  79.54759, 72.67453, 62.59805, 60.4373, 65.24623, 67.21675, 66.1386,
    62.37349, 61.10526, 56.61427, 46.86574, 47.47621, 49.14277, 49.91992,
    48.85139, 49.62273, 49.6862, 47.61465, 47.98009, 49.10149, 49.87043,
    50.41814, 50.59225, 52.56386, 52.65257, 44.65054, 38.40132, 37.20174,
    34.97364, 33.0242,
  85.46652, 81.4455, 76.75305, 76.08572, 78.23039, 76.58862, 76.59841,
    72.86924, 71.65776, 63.50576, 55.04935, 59.44603, 61.53169, 62.86357,
    60.56028, 59.10833, 57.40248, 54.18615, 51.31891, 51.10955, 51.00444,
    50.7317, 50.37095, 50.16636, 51.7122, 51.59298, 45.51232, 39.21423,
    37.2257, 34.23186,
  85.35552, 82.90147, 74.93615, 73.97845, 74.57152, 72.63066, 71.8637,
    73.7776, 77.18732, 68.99395, 61.0948, 65.48618, 67.37785, 68.38385,
    66.29863, 64.31525, 60.92505, 58.52291, 56.74409, 55.01093, 54.30135,
    53.1375, 50.53041, 48.82763, 50.08766, 52.75505, 52.16541, 44.53247,
    40.02811, 36.43105,
  92.34657, 89.99588, 85.36785, 78.13313, 75.532, 74.0686, 77.70721,
    80.77448, 76.98663, 68.5892, 67.43185, 69.37832, 70.18192, 67.8124,
    63.91632, 62.69605, 61.00448, 59.66058, 59.368, 57.91279, 56.74418,
    55.12051, 51.82924, 49.54239, 50.51883, 52.02907, 53.13142, 46.79454,
    38.15741, 35.60254,
  93.79298, 89.70723, 80.47741, 75.44266, 73.00391, 70.6013, 75.37184,
    75.5595, 69.58791, 64.84499, 67.37447, 68.73845, 69.23027, 67.5577,
    65.97144, 64.63875, 63.72063, 63.75607, 64.84459, 65.08354, 65.92336,
    67.55314, 66.29282, 62.84464, 62.17973, 62.64524, 63.74492, 56.30997,
    40.92905, 33.7893,
  93.7859, 86.62829, 82.23373, 80.24261, 80.34491, 77.30572, 76.27394,
    70.82508, 63.03663, 64.22789, 66.79096, 70.52257, 72.78986, 73.2489,
    73.65837, 72.12035, 70.10182, 70.54939, 73.29767, 74.68222, 71.55509,
    66.82281, 62.42377, 60.69723, 61.22379, 62.32705, 63.10211, 63.22641,
    54.4595, 38.02998,
  81.64459, 78.33313, 79.8802, 80.42173, 81.63239, 82.48114, 73.45258,
    62.54904, 58.68654, 61.188, 61.99037, 64.32614, 66.62209, 68.06138,
    68.98386, 68.73331, 66.53334, 64.08232, 60.5735, 56.741, 54.4379,
    52.23891, 48.86948, 46.73232, 47.64309, 48.81474, 48.46947, 46.21396,
    45.20625, 39.95474,
  80.42261, 80.52652, 77.57126, 74.90218, 78.60244, 86.06626, 86.20807,
    72.97482, 68.48816, 73.46603, 76.05322, 77.46423, 75.57506, 71.63643,
    66.70496, 61.55569, 53.74876, 46.98427, 45.34458, 43.85067, 42.02516,
    42.25903, 42.10212, 41.8022, 41.89546, 42.55177, 42.12627, 38.79184,
    35.51218, 32.9033,
  35.7547, 36.35471, 36.94776, 37.62001, 38.20327, 38.86774, 39.5541,
    40.27393, 41.00845, 42.05086, 43.7144, 44.0429, 42.13124, 42.81828,
    43.01071, 42.27581, 42.26202, 42.64497, 43.15816, 44.27591, 44.67594,
    43.62984, 44.27348, 46.55273, 48.47205, 48.20078, 50.34737, 51.01004,
    40.2493, 36.12956,
  39.86872, 40.89572, 41.02623, 42.39394, 42.64302, 43.06015, 44.09818,
    45.0533, 46.0675, 47.27238, 48.76246, 50.48141, 51.51149, 50.37695,
    49.70252, 49.99753, 49.02962, 49.57528, 50.50179, 51.34967, 51.34364,
    51.1472, 51.96483, 55.52448, 58.68625, 53.41549, 47.04934, 49.57439,
    40.80125, 37.17358,
  43.37062, 44.81845, 45.80369, 46.81992, 47.70693, 48.66246, 49.60611,
    50.72995, 51.99711, 53.16478, 54.37156, 55.93833, 57.32841, 58.89166,
    59.71132, 58.52628, 59.12689, 60.53744, 61.9867, 64.79593, 69.46017,
    73.5546, 73.28515, 70.73698, 68.31058, 63.10887, 55.67448, 48.15441,
    40.58832, 37.99646,
  50.36236, 52.03609, 53.61407, 55.22693, 56.38704, 57.50187, 57.59924,
    57.49538, 58.23681, 59.03734, 59.48888, 60.18333, 60.33728, 60.1498,
    62.61876, 64.01042, 62.13824, 60.96867, 64.41504, 68.68941, 74.40139,
    73.45755, 68.40443, 71.10561, 69.04277, 67.51112, 64.44337, 53.07123,
    42.21217, 36.81588,
  55.5126, 56.2087, 58.16493, 59.56639, 60.29695, 60.51464, 61.17043,
    61.87289, 63.57188, 64.43304, 64.48478, 66.42139, 67.36646, 67.49847,
    68.37913, 69.66187, 67.7543, 64.35409, 66.25098, 71.29561, 70.29246,
    61.44053, 61.671, 66.80428, 70.66689, 70.86327, 68.86004, 73.94518,
    67.08479, 44.53618,
  66.09026, 69.63686, 72.62254, 75.12121, 74.27667, 73.93773, 76.13129,
    76.51784, 76.56693, 78.11738, 81.63242, 89.9539, 96.87981, 93.31716,
    93.14117, 94.06113, 90.86255, 81.62578, 72.53828, 69.47594, 62.22541,
    54.84583, 59.25946, 62.88337, 66.8698, 67.06163, 67.59072, 78.64052,
    70.51767, 40.87915,
  72.85609, 76.18185, 78.95699, 81.45359, 81.84904, 84.3456, 90.80869,
    95.34019, 92.93663, 87.27347, 82.51019, 74.05013, 64.57408, 64.58867,
    65.44258, 67.16685, 67.15479, 62.96464, 57.8738, 58.26199, 56.00257,
    55.07214, 57.99938, 62.06791, 62.49277, 59.35325, 62.88947, 69.50603,
    58.00271, 34.77483,
  68.19917, 71.60074, 74.9919, 78.09056, 79.41678, 85.01173, 87.33591,
    73.65855, 66.27921, 66.36648, 63.78071, 61.01411, 58.99208, 59.22919,
    59.56747, 61.38083, 63.33504, 61.53194, 58.05414, 57.92602, 58.07294,
    59.88102, 62.97865, 64.54003, 62.2966, 62.57842, 68.50317, 67.35908,
    50.66625, 35.45062,
  77.36568, 80.5184, 82.86713, 84.31615, 85.87821, 87.37337, 80.10168,
    79.2701, 81.86641, 81.57784, 80.8201, 79.62997, 79.69076, 84.18684,
    85.09955, 76.46992, 74.93538, 75.19238, 73.02535, 67.88798, 65.8061,
    70.20487, 75.01917, 72.5495, 66.34141, 70.40955, 70.70635, 58.84175,
    38.41278, 35.87504,
  96.58352, 101.4828, 96.36072, 96.17589, 94.62751, 88.19922, 75.81868,
    81.59935, 81.53528, 83.27026, 85.07376, 86.96642, 84.46565, 81.5811,
    78.9286, 81.99618, 81.93388, 79.12868, 75.66241, 74.67228, 75.34222,
    72.82083, 68.7505, 63.10204, 66.69429, 73.52113, 65.44518, 44.38467,
    35.29649, 34.18799,
  115.3067, 114.9195, 114.3649, 101.3145, 103.0034, 92.34466, 84.4978,
    86.81107, 87.52155, 83.51665, 72.12913, 59.63668, 57.98799, 58.26662,
    59.09845, 60.56016, 62.07679, 62.27882, 62.72006, 65.1137, 70.45002,
    66.7298, 57.57487, 56.27109, 61.09017, 58.97774, 44.33688, 35.53488,
    35.75686, 34.26121,
  120.1843, 116.6631, 118.2098, 117.6621, 111.6129, 91.88791, 87.73718,
    80.42776, 74.2276, 68.72273, 64.08577, 60.9902, 62.80448, 62.45359,
    58.98911, 58.04311, 56.84239, 56.69202, 57.19458, 60.23949, 65.67277,
    63.96748, 57.35831, 63.42552, 65.32682, 51.33488, 36.91308, 39.27816,
    36.4718, 35.02169,
  126.5648, 126.5132, 126.503, 125.2648, 122.1994, 117.3719, 110.7047,
    101.563, 104.2054, 91.09584, 84.01007, 79.05558, 82.69717, 82.66611,
    73.60941, 61.43677, 62.04041, 60.80835, 59.89685, 62.35017, 63.81487,
    59.90955, 55.81855, 51.86396, 50.31177, 45.00667, 38.08176, 38.96206,
    38.06842, 35.94603,
  117.4722, 117.5646, 116.9685, 114.7337, 113.1714, 112.8266, 112.8331,
    111.7938, 108.891, 108.1026, 107.0683, 104.8318, 104.5432, 102.2177,
    91.07381, 76.14612, 70.335, 73.20197, 73.8092, 67.64045, 60.35922,
    53.81101, 48.16591, 41.95411, 38.41983, 38.05707, 36.79903, 36.13277,
    36.36563, 35.59451,
  94.82846, 90.57739, 91.3577, 91.70833, 92.35472, 95.03802, 100.4814,
    97.82626, 92.19025, 89.99509, 85.83562, 81.79882, 83.62227, 86.24442,
    84.48788, 80.43217, 73.12547, 68.3416, 66.68432, 61.71961, 50.82658,
    48.24464, 42.31145, 39.55362, 38.74234, 37.84292, 36.74294, 35.59182,
    34.94814, 34.56579,
  85.03383, 86.25876, 86.04201, 84.83209, 83.54495, 85.08332, 87.22507,
    82.39713, 75.88016, 72.26904, 70.87033, 67.65588, 66.4398, 70.71412,
    67.85822, 65.97405, 65.47636, 59.49215, 56.44704, 51.23969, 43.89934,
    44.0855, 40.41244, 39.29148, 38.80656, 37.768, 36.53528, 35.75753,
    35.06489, 34.55864,
  73.71729, 72.06835, 72.63428, 74.07697, 75.50897, 76.72334, 77.94099,
    78.79375, 77.09785, 73.26336, 68.97803, 74.22177, 79.34322, 74.07051,
    67.30342, 63.38863, 59.44582, 56.58566, 55.41731, 51.54834, 43.66928,
    44.09708, 41.14779, 39.2056, 38.41104, 37.94999, 36.22421, 34.89944,
    34.68676, 34.46841,
  67.56033, 68.34501, 67.61861, 69.43446, 71.18784, 73.20628, 74.83864,
    76.99324, 78.34559, 77.71765, 82.24126, 86.4099, 84.40873, 82.1505,
    76.97267, 69.81125, 64.61764, 62.80224, 62.32531, 55.48429, 45.05967,
    43.53569, 41.19529, 39.75695, 37.69928, 36.97002, 36.09124, 34.49261,
    34.37499, 34.2383,
  77.23466, 72.09093, 64.80897, 62.02404, 64.33194, 65.0223, 66.65161,
    68.37724, 68.78564, 70.75921, 74.0831, 72.27364, 67.74948, 69.88239,
    70.02149, 72.59753, 78.47444, 82.4268, 78.95353, 68.6474, 54.16426,
    46.52823, 42.5523, 40.57603, 38.17922, 36.86083, 35.98341, 34.7893,
    34.34128, 34.24663,
  75.86701, 70.5168, 62.48315, 57.92258, 59.19344, 59.5325, 60.40633,
    61.51987, 63.64348, 67.63498, 67.01442, 60.46403, 60.38478, 59.36295,
    58.06902, 58.31488, 62.16145, 67.50529, 68.59622, 66.15924, 59.89645,
    51.93549, 45.42204, 42.83287, 40.39116, 37.78919, 36.35149, 35.00074,
    34.32988, 34.26606,
  70.27576, 64.78025, 56.37395, 52.14329, 52.459, 52.86801, 53.85086,
    55.29137, 57.76797, 59.98866, 56.6741, 52.5882, 55.44794, 54.70539,
    52.78678, 51.74389, 52.81601, 54.53819, 56.15172, 56.05839, 55.91773,
    55.35993, 50.56118, 45.91505, 42.28846, 38.54877, 36.13373, 35.00933,
    34.36737, 34.29891,
  67.7048, 62.60875, 55.26922, 51.92918, 52.33569, 51.30397, 52.37461,
    53.45094, 56.58951, 56.93578, 51.37191, 48.91674, 50.77464, 50.56048,
    49.38594, 49.0026, 48.59854, 49.13505, 50.46597, 51.1259, 51.0191,
    50.49324, 50.68627, 49.51565, 45.19709, 39.52868, 36.73202, 35.69867,
    34.60079, 34.26179,
  71.00709, 69.36702, 61.17751, 58.62187, 61.08411, 61.41983, 60.07319,
    58.15904, 58.67736, 56.82066, 51.91999, 52.5255, 53.13326, 52.8828,
    51.40958, 51.10244, 50.11852, 48.20021, 47.8947, 47.93216, 47.58185,
    46.91196, 46.49313, 47.6957, 48.21791, 43.12119, 38.67725, 37.47383,
    35.82239, 34.40229,
  79.66855, 78.69725, 73.77067, 72.24744, 72.30078, 70.84458, 70.88467,
    70.50089, 72.25737, 68.11331, 63.20009, 65.28043, 65.86147, 65.55408,
    63.01495, 60.64255, 58.34085, 55.04388, 51.86744, 50.45817, 48.90395,
    47.57879, 46.67841, 46.44237, 47.76481, 47.76308, 43.66981, 39.29054,
    37.5168, 35.29304,
  81.82572, 77.59551, 70.79978, 68.72367, 68.81906, 67.7981, 68.42724,
    71.57621, 75.54497, 70.97182, 65.28296, 67.16039, 68.0414, 68.13869,
    66.13461, 64.0668, 60.68037, 57.7478, 55.33735, 52.92129, 51.28947,
    49.44118, 46.9985, 45.48201, 46.46646, 48.36228, 47.86896, 42.58953,
    39.18256, 36.64843,
  85.82576, 83.05438, 78.13908, 73.09121, 70.75835, 69.97279, 73.43626,
    77.76719, 76.83575, 71.49072, 70.40482, 70.93983, 71.03915, 69.24917,
    66.11613, 64.27169, 61.70871, 59.32962, 58.10007, 56.22952, 54.86765,
    53.35638, 50.29369, 47.86497, 47.75075, 48.25769, 48.5905, 43.80692,
    37.79828, 35.95267,
  86.86537, 84.30004, 78.19096, 74.70383, 72.47389, 70.64165, 74.26271,
    75.57823, 73.09094, 70.63492, 71.6333, 71.96394, 71.83986, 70.60536,
    68.36774, 66.24291, 64.12469, 62.54539, 61.86419, 60.60059, 60.11809,
    60.52366, 59.20341, 56.3036, 55.04452, 55.11519, 55.6769, 50.47513,
    39.93065, 34.98092,
  86.70231, 84.73213, 81.38506, 79.93347, 79.32564, 76.45747, 74.13794,
    70.08021, 65.36146, 65.21542, 65.77592, 66.76218, 67.40881, 66.92152,
    66.06509, 64.27303, 61.59862, 60.4571, 61.04258, 61.21307, 59.16961,
    56.06963, 53.28299, 52.1239, 52.44049, 53.2226, 53.72226, 54.24969,
    48.72087, 37.85169,
  72.68094, 72.04483, 72.83065, 73.02721, 74.17209, 75.56927, 69.51312,
    59.55502, 55.9977, 56.33298, 55.42369, 55.24409, 55.48814, 55.19951,
    54.86627, 54.40823, 52.74392, 51.18226, 49.44415, 47.77396, 46.91005,
    45.96632, 44.1886, 43.04607, 43.74375, 44.52301, 44.09311, 42.72306,
    42.46766, 38.79815,
  59.77789, 59.91107, 58.5611, 56.86637, 58.60056, 63.51352, 63.55066, 54.63,
    50.90057, 53.54527, 54.94926, 55.89648, 55.42957, 53.24221, 50.76431,
    48.94021, 44.81452, 41.33112, 40.83015, 40.19212, 39.2869, 39.61248,
    39.8128, 39.88518, 40.02285, 40.44168, 40.02442, 38.11722, 36.18069,
    34.39082,
  36.74014, 36.92252, 37.17819, 37.40199, 37.47905, 37.63744, 37.88586,
    38.21026, 38.57921, 39.24849, 40.43561, 40.37468, 38.52439, 39.08411,
    39.29816, 38.74894, 38.85566, 39.34613, 39.99028, 41.16376, 41.70905,
    40.96023, 41.64546, 43.63115, 45.4394, 45.81371, 48.14026, 49.22289,
    40.85547, 37.63162,
  39.59829, 39.97309, 39.77257, 40.40394, 40.07399, 39.93997, 40.34978,
    40.68699, 41.1051, 41.71201, 42.47329, 43.33103, 43.89887, 43.01985,
    42.55224, 43.09883, 42.61312, 43.57241, 44.84772, 45.99555, 46.33871,
    46.75099, 48.3047, 52.05605, 55.46391, 51.60682, 45.71345, 48.53208,
    41.20786, 38.43439,
  41.95002, 42.31183, 42.52582, 42.81578, 43.05658, 43.45318, 43.80799,
    44.26423, 44.842, 45.5053, 46.358, 47.60369, 48.91401, 50.39528,
    51.45163, 51.1719, 52.40539, 54.36346, 56.15049, 59.1496, 64.23094,
    69.60567, 70.25048, 66.65434, 63.51734, 59.28361, 53.29248, 47.42902,
    41.21195, 39.1886,
  47.68238, 48.65821, 49.69635, 50.88683, 51.91226, 52.95322, 52.90749,
    52.56775, 53.00807, 53.6894, 54.18308, 55.2179, 55.92087, 56.06419,
    58.73262, 60.59261, 59.36449, 58.78854, 62.05031, 65.92999, 71.81647,
    71.29143, 64.93311, 66.04139, 62.73962, 61.12164, 59.82554, 50.21923,
    41.40214, 38.00734,
  52.28141, 52.12629, 53.22915, 54.01656, 54.41586, 54.40064, 54.56522,
    54.68812, 55.5862, 56.04852, 56.02755, 57.43758, 58.66751, 59.52107,
    60.93599, 62.82503, 62.06273, 60.42285, 63.26064, 68.47964, 68.04117,
    58.79904, 57.81826, 61.65466, 64.35755, 64.59306, 63.15669, 68.00481,
    63.36139, 45.77866,
  57.51258, 59.71672, 61.94043, 64.17213, 64.05585, 64.44377, 67.35955,
    68.62143, 69.77522, 72.37225, 76.52689, 85.25107, 90.12112, 89.08664,
    88.60877, 88.2433, 86.67596, 82.04391, 73.8706, 70.54939, 62.99971,
    55.73079, 59.76073, 62.78753, 66.18617, 66.77502, 67.57255, 77.1535,
    69.8325, 42.24881,
  68.08565, 71.86224, 75.15646, 78.44574, 80.13435, 83.84799, 91.85768,
    92.5068, 91.51576, 90.77456, 87.51451, 79.68852, 70.98907, 70.71199,
    71.02522, 71.79824, 71.04109, 66.47354, 61.16212, 59.9171, 56.59539,
    55.33362, 58.21603, 61.87081, 62.61557, 60.57034, 64.41334, 70.40875,
    58.51931, 36.56408,
  69.70098, 72.702, 75.41553, 77.92999, 78.71658, 83.24947, 84.85308,
    71.15906, 63.12469, 61.95095, 58.49602, 55.20519, 53.21555, 53.79612,
    54.75444, 56.89551, 58.80643, 57.91822, 55.20967, 55.08736, 54.91333,
    56.33448, 59.69807, 62.22514, 61.50842, 62.98722, 69.73422, 68.22027,
    51.38997, 36.81376,
  71.69643, 72.89462, 73.90665, 74.26965, 75.06863, 74.91662, 65.84499,
    63.80484, 65.76682, 65.46159, 65.17142, 65.24962, 66.73282, 71.79294,
    73.43811, 66.89698, 67.12161, 68.69339, 67.47778, 63.59347, 62.30946,
    66.51564, 71.14785, 69.68714, 65.47456, 70.40578, 71.78275, 59.85647,
    39.90227, 37.49311,
  82.31203, 86.35895, 82.21567, 82.71738, 83.48183, 77.60387, 65.30374,
    71.35037, 72.41166, 75.01524, 78.03474, 81.89135, 80.70743, 78.53246,
    75.92554, 77.9396, 78.064, 76.14819, 73.94415, 73.25906, 73.93526,
    72.02782, 68.6452, 63.88078, 67.99432, 75.24992, 66.80974, 45.85323,
    36.79199, 36.21457,
  97.96635, 97.88544, 97.78906, 91.28238, 93.2521, 84.62299, 77.21396,
    81.10414, 82.72642, 80.00058, 71.38564, 60.85721, 59.89839, 60.16787,
    60.39732, 61.6352, 62.77815, 62.6461, 62.90198, 65.03326, 69.46938,
    66.22848, 58.40981, 57.13018, 62.01841, 60.4603, 46.50881, 36.97312,
    37.38582, 36.14693,
  101.4667, 98.34103, 100.2244, 99.71799, 97.99202, 81.85826, 79.55572,
    72.8253, 66.51688, 62.96098, 59.15171, 57.19628, 59.42481, 59.32732,
    56.83033, 56.50993, 55.95181, 56.06116, 56.42287, 58.84122, 63.85249,
    63.13454, 58.15084, 63.92881, 65.24385, 51.87421, 37.98135, 40.11398,
    37.95741, 36.8042,
  108.5335, 108.5943, 109.0323, 107.7838, 105.3697, 101.3483, 94.62504,
    80.8343, 86.79293, 76.25262, 71.28265, 68.41696, 72.65656, 73.6396,
    67.27623, 57.67076, 58.84302, 58.7612, 58.67019, 61.32915, 63.75655,
    61.7457, 58.73118, 55.13422, 52.3352, 46.21693, 39.51732, 40.52956,
    39.464, 37.64532,
  102.6823, 102.2346, 101.0886, 98.60837, 96.58242, 95.81357, 95.46661,
    94.78371, 92.76238, 92.53493, 92.61617, 90.82251, 90.53022, 90.28786,
    84.05578, 71.11972, 68.53259, 71.4929, 72.73589, 66.97096, 60.1502,
    55.32713, 50.87166, 44.1314, 40.47197, 39.96788, 38.73418, 38.05066,
    38.12818, 37.36121,
  90.5885, 86.17892, 87.2742, 86.88143, 87.61423, 90.01784, 94.00878,
    92.24799, 87.921, 87.82829, 84.17822, 79.84435, 81.10783, 81.93336,
    81.23813, 79.25672, 71.09736, 67.70616, 64.99721, 59.91635, 50.25077,
    48.00067, 42.6983, 40.34553, 39.98716, 39.38415, 38.45211, 37.4094,
    36.83312, 36.47837,
  78.7388, 80.75015, 80.95557, 80.09953, 78.76305, 79.60592, 80.83513,
    77.47615, 72.72321, 69.36868, 68.74004, 65.90556, 64.29022, 68.12299,
    65.39598, 63.25542, 63.18565, 57.89883, 54.75793, 50.13563, 43.65544,
    43.77808, 40.75078, 39.81589, 39.77079, 39.30694, 38.44307, 37.59333,
    36.8911, 36.48033,
  67.10172, 65.84178, 65.97176, 66.81295, 67.57484, 68.10351, 69.03893,
    70.33619, 69.14488, 66.11093, 62.16484, 66.29857, 70.80489, 66.74921,
    61.31729, 58.79538, 56.00444, 53.46716, 52.53521, 49.90979, 44.02921,
    44.17641, 41.48906, 39.93131, 39.68491, 39.54768, 38.1529, 36.93311,
    36.67304, 36.44464,
  62.23603, 62.96729, 62.06486, 63.14159, 63.95316, 65.1701, 66.43108,
    68.28793, 69.14957, 67.98238, 71.32712, 74.53923, 72.97699, 70.57971,
    65.08681, 60.20485, 56.06004, 55.35616, 55.7789, 51.81163, 44.65063,
    43.63922, 41.6835, 40.6227, 39.29504, 38.7467, 37.92287, 36.50367,
    36.3625, 36.2274,
  72.41509, 67.94607, 60.55398, 57.29439, 58.80631, 58.86079, 59.77101,
    60.87371, 60.76239, 62.37956, 65.5212, 64.19685, 59.87514, 61.05219,
    60.73041, 62.85364, 68.24245, 72.41518, 70.10358, 62.36271, 51.34576,
    45.66062, 42.73639, 41.28595, 39.55932, 38.55669, 37.75742, 36.68869,
    36.3184, 36.23757,
  69.83459, 65.61697, 58.46993, 54.53357, 55.99682, 56.50838, 57.25751,
    58.11158, 59.79499, 63.16457, 63.38577, 58.68014, 58.69723, 57.64873,
    56.41275, 56.81842, 60.00354, 64.24677, 64.53771, 61.87086, 56.33378,
    49.79952, 44.89425, 43.12587, 41.25313, 39.24694, 38.12306, 36.90975,
    36.32866, 36.26423,
  66.05473, 62.33441, 55.47075, 52.02251, 52.81754, 53.32816, 54.13708,
    55.08219, 56.85764, 58.85149, 56.51208, 53.07445, 55.31496, 54.57502,
    52.79731, 51.98779, 52.90438, 54.21188, 55.05596, 54.20956, 53.3828,
    52.4976, 48.82372, 45.53797, 42.73088, 39.92898, 37.96767, 36.93094,
    36.38201, 36.29243,
  63.84231, 60.59388, 54.19201, 51.27444, 51.66285, 50.85165, 51.62106,
    52.2858, 54.55851, 54.84615, 50.57159, 48.42185, 49.94249, 49.76015,
    49.04375, 48.95076, 48.83399, 49.25617, 50.14052, 50.42942, 50.11346,
    49.49674, 49.34233, 48.08201, 44.53908, 40.30739, 38.23368, 37.30529,
    36.4901, 36.26598,
  65.30231, 63.67616, 56.29307, 53.70573, 55.44678, 55.42733, 54.2219,
    52.4769, 52.8546, 51.22799, 47.16193, 47.66091, 48.4487, 48.92576,
    48.57027, 48.81269, 48.3715, 47.25172, 47.20564, 47.19889, 47.04501,
    46.54868, 45.83688, 46.29722, 46.21876, 42.35236, 39.2244, 38.46082,
    37.29177, 36.3371,
  72.41217, 71.90134, 66.63358, 64.7648, 64.44009, 62.94293, 62.61187,
    61.63544, 63.24108, 60.12407, 56.21222, 57.80332, 58.66341, 59.04313,
    57.56033, 56.08244, 54.51363, 52.11221, 49.67485, 48.59042, 47.76699,
    46.81531, 45.85995, 45.45038, 46.32699, 46.2092, 42.95985, 39.6303,
    38.40446, 36.91545,
  74.74477, 70.60573, 64.83658, 62.5567, 62.11723, 60.96293, 61.6493,
    64.36436, 67.93858, 64.04642, 59.69796, 61.48011, 62.69062, 63.38094,
    61.89819, 60.48549, 58.59775, 56.41505, 53.67638, 51.76261, 50.77155,
    49.21842, 46.91098, 45.68882, 46.63654, 48.06787, 47.19987, 42.75497,
    40.01791, 38.05263,
  78.55702, 75.19055, 69.64556, 64.95172, 62.88803, 61.99201, 64.88768,
    68.9448, 68.38438, 63.506, 62.83623, 63.79583, 64.54743, 63.6527,
    61.29631, 60.11444, 58.97846, 57.26662, 55.41239, 53.70158, 53.00328,
    51.51946, 48.25997, 46.44825, 46.74892, 47.06542, 47.17326, 43.66434,
    39.12975, 37.56526,
  80.38359, 75.87429, 70.03771, 65.98402, 63.9422, 62.28125, 65.3611,
    66.82509, 65.24766, 62.96578, 64.11939, 64.87588, 65.27614, 64.41516,
    62.69022, 61.16172, 60.36413, 59.73245, 58.43336, 57.3115, 57.66995,
    57.93346, 55.71147, 52.59172, 51.42163, 51.26099, 51.53392, 47.78541,
    40.17079, 36.74781,
  78.35177, 75.50745, 72.23322, 71.14268, 71.11115, 69.51479, 68.63452,
    66.32236, 63.38841, 63.77359, 64.93883, 66.24838, 67.20088, 67.15833,
    66.55513, 65.14922, 63.55915, 62.86263, 62.53856, 62.0829, 60.69202,
    57.9711, 54.41331, 52.33128, 51.99122, 52.1339, 52.2384, 52.41363,
    47.45547, 38.88988,
  65.34229, 65.24962, 65.99393, 66.46956, 68.50111, 70.64552, 66.85826,
    59.42046, 56.76816, 57.49818, 57.42867, 58.02468, 58.9527, 59.43171,
    59.59432, 59.3463, 58.24496, 56.88853, 54.66383, 52.53203, 51.2742,
    49.89514, 47.76466, 46.17075, 46.08167, 46.13509, 45.57322, 44.39335,
    43.74585, 40.22134,
  59.08384, 59.72306, 59.54836, 59.13517, 61.48935, 66.42888, 66.64801,
    58.82108, 55.27443, 57.44632, 58.93211, 60.07833, 59.64399, 57.44262,
    54.82862, 52.75383, 49.18119, 46.44816, 45.71276, 44.64128, 43.58113,
    43.56453, 43.36283, 42.97876, 42.60398, 42.28085, 41.46963, 39.9817,
    38.2904, 36.51377,
  39.97648, 39.99686, 40.07787, 40.08947, 40.10538, 40.18114, 40.31079,
    40.57906, 40.87459, 41.37465, 42.25691, 42.07695, 40.60912, 40.93608,
    41.10846, 40.71003, 40.64118, 40.79262, 40.99904, 41.64562, 41.94559,
    41.28806, 41.55728, 42.90143, 44.36596, 44.91094, 46.89195, 48.43936,
    43.25467, 40.95912,
  40.92988, 41.0479, 40.82217, 41.1926, 40.95164, 40.89402, 41.21799,
    41.5632, 41.93567, 42.37847, 42.87886, 43.25536, 43.28294, 42.47032,
    41.97615, 42.16818, 41.46991, 41.74767, 42.3567, 42.93324, 43.06951,
    43.48484, 45.51353, 50.0898, 54.29351, 51.35571, 46.68608, 49.31486,
    43.72438, 41.52195,
  40.59973, 40.52532, 40.50914, 40.51706, 40.51332, 40.70146, 40.87546,
    41.10229, 41.42787, 41.71528, 42.01495, 42.51765, 43.00823, 43.59024,
    44.00785, 43.62215, 44.40776, 45.85967, 47.29673, 50.28296, 55.63943,
    62.13631, 64.97375, 64.05008, 62.48474, 57.87935, 53.51735, 48.77787,
    43.89843, 42.26961,
  40.74085, 41.04906, 41.78537, 42.60277, 43.32657, 44.18941, 44.36047,
    44.21984, 44.61648, 45.24639, 45.50423, 46.102, 46.60042, 47.02002,
    49.50546, 51.66072, 52.07072, 52.96231, 57.07812, 62.63884, 70.05343,
    70.84738, 65.22818, 65.53239, 62.09048, 60.24296, 58.75945, 50.52368,
    43.34405, 41.17543,
  43.53876, 43.55465, 44.70536, 45.61044, 46.10678, 46.13659, 46.01818,
    45.8409, 46.28112, 46.30962, 45.87582, 46.63593, 47.95208, 49.94335,
    52.67064, 55.92039, 57.46648, 58.15278, 62.31398, 67.93162, 68.02066,
    59.35622, 56.63801, 59.78969, 61.58813, 61.29093, 60.62794, 65.51809,
    62.93895, 48.52127,
  44.84528, 45.65121, 46.96633, 48.09628, 47.29543, 46.33961, 47.35607,
    48.26321, 50.06517, 53.51757, 58.80139, 68.65953, 77.66357, 77.28407,
    80.00649, 81.74472, 81.14178, 77.62029, 71.61669, 68.57642, 61.32587,
    53.73783, 57.74022, 61.29015, 65.50059, 67.19287, 69.21954, 78.41093,
    73.80611, 46.269,
  47.67075, 49.87206, 52.55666, 55.55465, 58.0188, 62.78481, 72.00587,
    81.01396, 81.8082, 81.8619, 81.93499, 81.66082, 75.48167, 75.52504,
    75.98967, 76.44646, 76.11402, 70.80336, 64.17435, 62.00524, 58.24188,
    57.36283, 60.89303, 64.70805, 66.48079, 65.49005, 69.39902, 75.35712,
    62.68452, 40.15692,
  57.61029, 62.44007, 67.25085, 72.55636, 77.09352, 82.41881, 83.10514,
    81.161, 74.62239, 73.17455, 68.80812, 63.80167, 60.22388, 59.74986,
    59.81945, 61.35186, 62.50938, 60.76473, 57.9167, 57.70943, 57.32529,
    58.43441, 61.22224, 63.43796, 62.92883, 64.09152, 69.87171, 69.01257,
    54.49773, 40.13068,
  69.159, 73.04066, 75.77091, 77.65012, 79.69707, 79.45622, 69.28767,
    63.85157, 62.98229, 61.04129, 59.29228, 58.36412, 59.14352, 63.37897,
    65.73038, 61.85497, 63.00031, 65.18549, 64.58967, 61.45657, 60.50929,
    64.3025, 68.69077, 68.16661, 66.13789, 72.17297, 74.60858, 63.37915,
    43.63005, 40.82528,
  76.16846, 79.52161, 75.88789, 75.70779, 75.63828, 69.12287, 55.40489,
    59.55229, 60.52538, 63.64448, 67.66152, 71.46624, 71.20456, 70.50967,
    69.3232, 71.75658, 73.6078, 73.49346, 72.18593, 71.43748, 72.59717,
    72.04423, 69.93386, 66.38843, 70.6293, 78.11012, 70.78403, 49.89584,
    40.18802, 40.02844,
  75.82093, 75.68953, 75.28737, 74.11073, 76.91994, 71.3703, 65.77348,
    71.73592, 76.45053, 77.7376, 71.83185, 62.91981, 61.33736, 61.85044,
    62.81908, 64.53162, 66.00117, 66.39748, 66.96701, 68.88826, 72.72691,
    69.99866, 63.60307, 62.68208, 67.65626, 65.90201, 51.39485, 40.47613,
    40.72972, 39.88916,
  80.84531, 75.05933, 81.84559, 86.81628, 83.58121, 75.1729, 77.56979,
    72.39767, 67.06953, 65.41995, 60.80017, 57.8927, 60.0421, 60.6813,
    59.64251, 60.34706, 59.9077, 60.18972, 60.45572, 62.34039, 66.49024,
    65.61012, 61.39244, 66.46367, 67.76199, 55.2622, 40.99467, 42.62167,
    41.36385, 40.38984,
  90.76937, 93.04118, 95.40824, 95.50797, 93.99507, 90.66337, 83.96831,
    71.3998, 76.54578, 68.758, 65.18858, 63.79914, 68.1611, 70.0566,
    65.79258, 57.71545, 59.27108, 59.35477, 59.7971, 62.63651, 65.84212,
    65.32696, 63.03468, 59.32321, 55.86283, 49.21469, 42.22742, 43.68016,
    42.60615, 41.1391,
  94.46458, 95.5779, 94.53082, 91.30999, 88.40197, 86.27757, 85.00987,
    84.48754, 82.89273, 82.79784, 83.06931, 82.04068, 82.26514, 82.30007,
    78.46384, 68.63101, 67.24473, 72.19408, 74.50283, 70.41747, 65.56464,
    60.93711, 55.501, 48.887, 44.91601, 43.85281, 42.49428, 41.93872,
    41.74769, 40.98263,
  89.94793, 88.61542, 86.6162, 84.5882, 83.44161, 84.26665, 86.37983,
    85.9865, 84.12727, 83.65388, 82.84697, 79.62019, 79.58492, 81.85091,
    81.20327, 80.22624, 76.52143, 73.32407, 70.99133, 65.50461, 55.56861,
    52.04569, 46.38261, 43.49479, 43.16629, 42.81698, 42.03455, 41.10303,
    40.60722, 40.2369,
  84.48949, 84.07306, 84.14317, 83.11543, 82.32828, 83.38835, 84.36914,
    81.18312, 76.58922, 73.01849, 72.00126, 69.81673, 70.02906, 73.4714,
    71.01139, 69.4666, 68.27137, 62.64753, 58.84017, 53.72321, 47.44394,
    46.58214, 43.4398, 42.64708, 42.7905, 42.4801, 41.78162, 41.02427,
    40.44922, 40.13766,
  75.63802, 74.00809, 73.06784, 72.43416, 71.66856, 70.64229, 70.41797,
    70.95168, 69.53278, 66.8932, 63.64933, 66.71692, 70.72724, 67.86671,
    63.14824, 60.40907, 57.64947, 54.93511, 54.00728, 51.37233, 46.40336,
    46.5814, 44.0284, 42.72568, 42.60356, 42.5642, 41.57512, 40.61601,
    40.33736, 40.13001,
  64.79489, 64.50677, 63.43143, 63.61689, 63.76993, 64.38252, 65.10281,
    66.4842, 67.01267, 65.85859, 68.11108, 70.78579, 69.51896, 67.24082,
    62.87374, 58.60429, 54.33608, 53.37203, 54.26223, 51.67351, 46.55898,
    46.13056, 44.31231, 43.3801, 42.43329, 42.00356, 41.31078, 40.23928,
    40.11648, 39.98009,
  70.21181, 66.80715, 60.65702, 57.71447, 59.03797, 59.0153, 59.60223,
    60.24154, 59.8784, 60.85608, 63.14272, 61.49416, 56.76727, 56.66098,
    55.68082, 56.71021, 61.17043, 65.64498, 65.29233, 60.06113, 51.92425,
    47.47372, 44.98014, 43.94846, 42.54837, 41.75125, 41.09775, 40.27784,
    40.03976, 39.95341,
  69.80554, 65.11477, 57.91151, 53.83524, 54.63947, 54.39332, 54.50484,
    54.77402, 55.85227, 58.6203, 58.94123, 55.05376, 55.003, 54.75826,
    54.69926, 56.17163, 60.0382, 64.32706, 64.40834, 61.24397, 55.79655,
    50.1422, 46.20275, 45.18822, 43.76065, 42.3404, 41.39877, 40.44818,
    40.02093, 39.96338,
  66.5295, 62.74504, 55.4268, 51.65778, 52.14722, 52.26875, 52.791, 53.71959,
    55.6799, 57.9333, 56.51127, 54.30271, 56.92135, 56.94658, 56.02964,
    55.75426, 56.47802, 56.93399, 56.52474, 54.68045, 53.27706, 52.14485,
    49.32444, 47.13406, 45.23112, 43.18597, 41.48944, 40.53231, 40.08168,
    39.98071,
  64.31178, 61.44627, 55.19046, 52.26937, 52.80958, 52.56993, 53.79323,
    54.89172, 57.25787, 57.78437, 54.48363, 52.93354, 54.20223, 53.78896,
    52.82076, 52.30402, 51.60278, 51.22913, 51.39476, 51.46541, 51.46329,
    51.11448, 50.80944, 49.61636, 46.90649, 43.39575, 41.63509, 40.83073,
    40.14478, 39.99074,
  63.36525, 61.86362, 55.2719, 53.05312, 55.00765, 55.58035, 55.37725,
    54.36977, 54.61066, 53.04912, 49.35435, 49.49369, 49.99736, 50.02905,
    49.56051, 49.89624, 49.87488, 49.17273, 49.23074, 49.37363, 49.42614,
    49.12173, 48.39828, 48.2367, 47.71399, 44.37427, 42.11765, 41.55493,
    40.69845, 40.04319,
  65.85736, 65.35512, 60.56075, 59.26654, 59.62592, 58.54527, 58.21851,
    57.38508, 58.36916, 55.58397, 52.29715, 54.15138, 55.45326, 56.2171,
    55.54844, 55.22014, 54.57359, 53.02079, 50.9682, 49.8265, 49.35122,
    48.88224, 47.90869, 47.34212, 47.69825, 47.20137, 44.7983, 42.38937,
    41.50145, 40.47491,
  68.02027, 65.11215, 59.48172, 57.23126, 56.98032, 55.90619, 56.37642,
    58.64071, 62.03175, 59.27678, 56.06376, 58.34069, 60.09706, 61.122,
    60.38012, 59.78578, 58.74311, 57.09627, 54.5333, 52.82362, 52.11335,
    50.86685, 48.82212, 47.66305, 48.25992, 49.20023, 48.40842, 44.8788,
    42.90251, 41.45131,
  70.07996, 68.22325, 62.48094, 58.05201, 56.86478, 56.46699, 59.32716,
    63.60202, 64.33646, 60.4315, 60.1282, 61.67207, 62.85421, 62.3756,
    60.60828, 60.13447, 59.75501, 58.47204, 56.64391, 55.19078, 54.31393,
    52.69271, 49.88027, 48.42974, 48.79363, 48.86906, 48.77809, 45.98663,
    42.44232, 41.12639,
  71.25336, 68.18852, 62.62379, 58.86298, 57.71921, 56.99833, 60.10059,
    62.37521, 61.86539, 59.95836, 61.20842, 62.0919, 62.41573, 61.73451,
    60.53798, 59.6667, 59.36982, 58.98161, 58.02267, 57.15543, 57.04498,
    56.83959, 55.12863, 53.12446, 52.50761, 52.06699, 51.95729, 48.7679,
    42.82556, 40.37055,
  71.23396, 67.65057, 64.11554, 63.05418, 63.49214, 62.75776, 62.76636,
    61.78175, 59.93088, 60.08894, 61.18022, 62.217, 62.96317, 63.17232,
    63.14758, 62.69011, 62.28078, 62.18681, 62.29565, 62.42567, 60.98637,
    58.3668, 55.56385, 54.01621, 53.67456, 53.32513, 52.53071, 51.90799,
    48.19154, 41.92041,
  63.11615, 62.31941, 62.72908, 63.21066, 65.25382, 67.3962, 64.85301,
    59.43649, 57.78208, 58.37519, 58.44823, 59.10874, 60.22613, 61.58567,
    62.6605, 63.04031, 62.59765, 61.64775, 59.67339, 57.52072, 55.66964,
    53.85896, 52.03149, 50.68443, 50.47048, 50.02551, 48.95456, 47.35077,
    46.08725, 43.08062,
  59.14109, 59.55077, 59.73058, 59.60169, 61.69809, 66.09024, 66.43826,
    60.24446, 57.64065, 59.24766, 60.39016, 61.3608, 61.47018, 60.41293,
    59.03708, 57.53083, 54.85852, 52.48026, 51.2658, 49.72645, 48.31403,
    47.97091, 47.71732, 47.34754, 46.86707, 46.34805, 45.27033, 43.59103,
    42.13137, 40.46934,
  39.4051, 39.34304, 39.371, 39.38811, 39.38274, 39.42865, 39.48822,
    39.63077, 39.82029, 40.14752, 40.76317, 40.71166, 39.6337, 39.82361,
    39.95384, 39.74654, 39.76357, 39.86563, 39.99321, 40.49039, 40.71047,
    40.0326, 40.03303, 40.8584, 42.02, 42.62604, 44.03077, 45.72609,
    41.86938, 40.1566,
  39.99566, 40.0572, 39.86048, 40.08928, 39.87093, 39.76209, 39.99865,
    40.2701, 40.60376, 40.99529, 41.38316, 41.55579, 41.50475, 40.98987,
    40.63724, 40.9142, 40.45819, 40.60493, 40.89095, 40.95959, 40.39925,
    40.07804, 41.73159, 46.35571, 51.08604, 48.87418, 44.28502, 47.13831,
    42.57125, 40.7201,
  40.10006, 40.0673, 39.9896, 39.92921, 39.80764, 39.88062, 40.02869,
    40.24408, 40.44277, 40.60115, 40.79631, 41.117, 41.35337, 41.58607,
    41.71737, 41.09036, 41.14326, 41.55235, 41.70283, 43.34245, 47.89409,
    54.98154, 59.45909, 60.19664, 59.55264, 54.99379, 51.15492, 46.79177,
    42.76583, 41.41137,
  40.1399, 40.1839, 40.50002, 40.9183, 41.23054, 41.76952, 41.90223,
    41.78253, 42.11513, 42.62342, 42.82034, 43.20509, 43.29167, 42.91714,
    43.935, 44.78744, 44.45458, 44.58997, 48.18407, 54.55942, 63.95788,
    67.42642, 62.63237, 62.56253, 59.18816, 57.80094, 56.51067, 48.24535,
    41.79617, 40.23446,
  41.05016, 40.91058, 41.77874, 42.65269, 43.42602, 43.82531, 44.05313,
    43.90006, 43.88378, 43.23705, 41.8186, 41.06971, 40.82368, 41.55946,
    43.2065, 45.82272, 48.07116, 50.79681, 57.45291, 65.40779, 67.55843,
    59.49641, 54.82702, 57.08454, 57.81345, 57.27542, 56.23656, 60.90864,
    60.13425, 47.91732,
  42.11873, 43.005, 44.25554, 45.19598, 44.28926, 42.70013, 41.91892,
    40.86728, 40.50765, 41.64198, 45.19093, 53.54829, 62.74104, 63.51924,
    68.15903, 73.28072, 74.19753, 73.46392, 71.97601, 69.21831, 60.30607,
    50.23083, 53.03005, 55.81697, 59.3237, 60.99795, 63.15227, 71.80589,
    71.43732, 46.6538,
  42.972, 43.56296, 44.1358, 44.48573, 44.15729, 45.60815, 52.12547,
    61.54568, 66.51553, 69.38582, 73.15767, 72.81071, 69.6997, 72.56765,
    75.70913, 75.89078, 75.54294, 72.70846, 64.53822, 59.87529, 53.87879,
    51.93213, 56.02373, 60.05947, 62.86948, 63.26932, 67.93483, 72.2535,
    62.66116, 39.66109,
  43.05856, 44.48113, 47.17431, 51.11688, 55.9814, 66.48439, 75.94391,
    72.84187, 69.89229, 71.68165, 69.97727, 66.58206, 64.41756, 64.99799,
    64.60254, 64.44164, 63.11226, 58.95725, 54.58358, 53.74705, 53.54865,
    55.32401, 58.81341, 61.91724, 62.36113, 63.7887, 69.73027, 69.14626,
    54.06755, 39.42673,
  48.75022, 53.21904, 58.5675, 64.33499, 71.7652, 76.27625, 70.62085,
    66.01357, 65.93934, 64.5015, 62.39129, 61.00095, 61.03218, 63.13981,
    63.4116, 58.7375, 58.02543, 59.04694, 58.83664, 57.01743, 56.98089,
    60.66064, 64.80059, 65.28877, 64.23511, 70.57393, 73.21363, 64.0633,
    42.99308, 39.95097,
  62.31121, 69.46968, 70.08085, 74.08598, 77.59902, 73.88198, 58.17641,
    60.89872, 60.69815, 62.31314, 64.8138, 67.39581, 66.94571, 65.68001,
    63.40255, 64.2637, 65.92423, 66.26715, 65.65674, 65.49603, 67.25881,
    67.81681, 66.5578, 63.41763, 66.98556, 73.62112, 71.85033, 50.51442,
    39.52883, 39.486,
  71.28663, 75.78828, 76.1356, 74.43347, 76.01366, 67.74037, 59.57567,
    65.54272, 70.00001, 72.50032, 68.36678, 60.8698, 59.06597, 58.81028,
    58.9, 60.67557, 62.16275, 62.67222, 63.6118, 65.9054, 70.02611, 68.57167,
    62.86526, 62.33124, 68.10823, 67.99501, 53.40011, 39.98079, 40.01267,
    39.28918,
  77.3074, 69.49499, 71.91051, 74.68716, 72.57569, 66.22434, 72.43061,
    69.92735, 64.91861, 64.6504, 59.2835, 55.27914, 57.34081, 58.09336,
    57.24967, 58.59106, 58.66629, 59.26918, 59.76415, 61.68302, 65.7364,
    65.4198, 61.73725, 66.56306, 68.23766, 56.55293, 40.49167, 41.43131,
    40.53269, 39.67154,
  80.12678, 81.46468, 85.09438, 87.42754, 88.17151, 86.77541, 80.9029,
    65.91573, 70.79839, 64.05972, 59.95498, 60.02852, 65.33444, 67.74934,
    64.41126, 56.36073, 57.66541, 58.03115, 58.58105, 61.36709, 65.4549,
    66.59877, 65.08956, 61.19085, 56.23744, 48.65128, 40.91077, 42.72233,
    41.49393, 40.40094,
  85.06134, 89.33416, 91.38106, 89.84419, 87.18279, 83.64766, 80.35247,
    79.49452, 76.68726, 77.31746, 78.82635, 77.71305, 77.81684, 77.61544,
    74.54901, 63.93445, 63.22768, 68.70647, 72.76366, 70.62301, 67.86183,
    63.44781, 56.89484, 49.68737, 44.78312, 43.10829, 41.77657, 41.32103,
    40.91145, 40.30241,
  88.4128, 89.4221, 86.76342, 83.24157, 80.07128, 79.47548, 81.52493,
    81.98345, 80.32765, 80.14436, 79.44039, 78.05534, 76.8327, 77.23539,
    76.24702, 74.93463, 73.84158, 73.93295, 73.5138, 68.53122, 58.46098,
    53.37681, 46.53321, 42.77567, 42.45994, 42.15181, 41.36328, 40.48804,
    40.01919, 39.64499,
  85.72818, 84.06142, 81.87624, 79.97672, 79.36359, 80.63452, 81.94427,
    81.40327, 78.34583, 74.30121, 71.89458, 69.13445, 69.8006, 74.21119,
    73.36455, 72.39916, 71.4389, 66.23979, 61.43099, 55.01645, 47.90164,
    45.78317, 42.41425, 41.69284, 42.04671, 41.82206, 41.01969, 40.32887,
    39.80611, 39.53125,
  80.92261, 77.46765, 76.92865, 77.27931, 77.36205, 75.92905, 74.15602,
    73.19638, 70.48228, 67.36344, 65.04713, 68.17525, 72.65355, 71.27078,
    66.67047, 63.3841, 59.63577, 55.41454, 52.82351, 49.66547, 44.96098,
    44.79998, 42.66579, 41.63946, 41.67719, 41.68468, 40.83178, 39.99733,
    39.69291, 39.52616,
  72.23116, 72.54305, 71.98824, 71.35399, 69.67809, 68.28372, 67.66777,
    68.13728, 68.36088, 67.72793, 70.25002, 73.15755, 72.26804, 69.101,
    63.32346, 58.41995, 53.20397, 50.53258, 50.51041, 48.43721, 44.47761,
    44.49484, 42.9335, 42.1182, 41.53649, 41.19743, 40.58423, 39.69261,
    39.52837, 39.39959,
  77.64977, 75.11021, 68.74474, 64.42931, 64.66543, 64.34647, 65.00193,
    65.95913, 65.99812, 66.94319, 68.61842, 66.2094, 60.06913, 57.39377,
    53.75451, 52.56753, 54.6907, 57.69867, 58.14691, 55.07647, 49.36834,
    45.89863, 43.5517, 42.83962, 41.69023, 41.08453, 40.48552, 39.67065,
    39.44492, 39.36129,
  78.39842, 72.96919, 65.40263, 61.11933, 62.29048, 62.34919, 62.51505,
    62.4528, 62.2814, 62.86191, 61.24294, 55.75007, 53.23326, 51.18939,
    49.81912, 50.83018, 54.56913, 59.20507, 60.17756, 57.7621, 53.10832,
    48.07525, 44.55043, 43.92274, 42.76198, 41.56025, 40.73642, 39.85877,
    39.39394, 39.37977,
  74.32687, 69.98424, 62.89376, 58.98125, 59.38799, 58.73663, 58.03114,
    57.29033, 56.99514, 56.7388, 53.9186, 51.06601, 52.74061, 52.89341,
    52.82748, 53.78965, 55.53685, 56.46983, 55.57029, 52.7471, 50.52414,
    49.05854, 46.9442, 45.43858, 43.99569, 42.35389, 40.89772, 39.95924,
    39.43917, 39.38854,
  70.85316, 67.46896, 60.59799, 56.42477, 55.95518, 54.42162, 54.1342,
    53.97541, 55.047, 55.10049, 52.50596, 51.95354, 54.05213, 54.56346,
    54.35994, 54.04076, 52.98876, 51.6839, 50.56353, 49.49014, 48.91909,
    48.74345, 48.75336, 47.40099, 45.2872, 42.61559, 41.07042, 40.21662,
    39.53357, 39.40751,
  67.86368, 65.08318, 57.43753, 53.69419, 54.68542, 54.48338, 54.15764,
    53.68464, 54.33508, 53.82583, 51.63187, 52.29827, 53.06546, 52.85608,
    51.73036, 50.91864, 49.77236, 48.45358, 48.11894, 48.04284, 48.04334,
    47.88288, 47.34482, 46.46813, 45.81282, 43.15032, 41.24643, 40.73638,
    39.99805, 39.47056,
  67.4221, 65.95249, 60.34107, 58.17522, 58.3982, 57.48009, 57.36911,
    56.97979, 58.3236, 56.88577, 54.50581, 55.71543, 56.44609, 56.13686,
    54.52946, 53.53554, 52.6595, 51.49257, 49.85881, 48.79358, 48.22629,
    47.77036, 46.72683, 45.69192, 45.72446, 45.27095, 43.41446, 41.49174,
    40.71665, 39.80914,
  69.52982, 66.95674, 60.82557, 58.07822, 57.63717, 56.43496, 57.01054,
    59.03164, 61.97567, 59.67086, 56.83985, 58.21206, 59.24397, 59.45149,
    58.26048, 57.66213, 56.76386, 55.36734, 53.0234, 51.3269, 50.46442,
    49.27451, 47.23331, 46.07842, 46.56348, 47.04031, 46.13228, 43.26983,
    41.77999, 40.63617,
  70.55832, 68.44157, 62.61575, 58.37959, 57.27788, 56.63887, 59.12445,
    63.05337, 63.88836, 60.21301, 59.61881, 60.83202, 61.92609, 61.44263,
    59.58829, 59.15386, 58.56985, 57.12628, 55.10708, 53.50362, 52.28747,
    50.54371, 48.02095, 46.98133, 47.42062, 47.16464, 46.82813, 44.49411,
    41.63673, 40.49492,
  70.74598, 68.0626, 62.39705, 58.7569, 58.20296, 57.52576, 60.1255,
    62.35273, 62.16838, 60.25919, 61.21173, 61.97588, 62.42197, 61.31771,
    59.57459, 58.78189, 58.05031, 56.8708, 55.28688, 54.18866, 53.73725,
    53.36111, 52.11085, 50.66108, 50.07475, 49.36032, 49.10358, 46.69323,
    41.85836, 39.79548,
  70.36565, 67.08993, 63.2502, 61.82249, 62.8149, 62.53235, 62.98132,
    62.71786, 61.15688, 61.1305, 61.82915, 62.27344, 62.64729, 61.92224,
    60.74941, 59.94877, 59.21455, 58.55613, 58.56649, 58.99424, 58.03401,
    55.87442, 53.20341, 51.56108, 50.99684, 50.33795, 49.65432, 48.94447,
    45.80403, 40.93973,
  63.19803, 62.4496, 62.57405, 62.78997, 64.60391, 66.7493, 65.11695,
    60.70593, 58.90698, 59.12695, 58.76749, 58.99879, 59.75838, 60.36977,
    60.67761, 60.87245, 60.51277, 59.72144, 58.34724, 56.76006, 54.95712,
    53.01997, 51.08295, 49.59779, 49.22594, 48.73593, 47.85037, 46.28153,
    44.68675, 41.99407,
  59.16629, 59.70018, 59.9986, 59.68581, 61.35391, 65.07019, 65.66043,
    60.22798, 57.65334, 58.53241, 59.13901, 60.10423, 60.52687, 59.75208,
    58.68256, 57.70726, 55.46002, 53.23051, 51.94793, 50.18721, 48.5901,
    48.03902, 47.65703, 47.15971, 46.63153, 45.9279, 44.70567, 43.01796,
    41.5395, 39.99693,
  6.25687, 5.190001, 5.619899, 5.682805, 5.771177, 5.889614, 6.105238,
    6.380556, 6.839632, 7.774556, 8.712325, 10.1572, 12.05477, 15.01349,
    18.32574, 22.38458, 26.88154, 32.11287, 38.09879, 44.5669, 51.10794,
    56.55153, 60.58245, 63.12096, 64.29952, 64.35441, 64.48012, 64.84978,
    63.78711, 62.12142,
  4.52338, 3.710723, 4.102583, 4.218025, 4.289217, 4.315365, 4.398911,
    4.466805, 4.609581, 5.009672, 5.943151, 7.628005, 10.14161, 13.12553,
    16.86249, 21.29286, 26.55811, 32.54815, 38.9595, 45.99526, 52.23207,
    57.73803, 61.7994, 64.29839, 65.31686, 64.79241, 64.06286, 64.57356,
    63.88699, 62.61365,
  6.089709, 4.957926, 5.406588, 5.371065, 5.528627, 5.645888, 5.756649,
    5.855119, 6.032568, 6.445126, 7.348707, 8.99094, 11.4396, 14.60743,
    18.2303, 22.42577, 27.52895, 33.53497, 40.35846, 47.69859, 54.6811,
    60.20358, 64.02855, 65.84795, 66.15834, 65.66779, 65.2196, 64.36484,
    63.47738, 62.5569,
  6.028405, 4.87332, 5.318094, 5.28399, 5.440973, 5.587934, 5.728473,
    5.875947, 6.233828, 6.966797, 8.241919, 9.996846, 12.28163, 15.42115,
    19.30611, 23.53521, 28.41892, 33.69344, 40.27237, 47.67628, 54.95227,
    60.61676, 63.88735, 66.02084, 66.40971, 66.47053, 66.53735, 65.56525,
    64.35278, 63.40775,
  6.48675, 5.361508, 5.837393, 5.78323, 5.865902, 5.859488, 5.926966,
    6.008107, 6.411301, 7.369625, 8.936207, 11.17256, 13.77176, 16.95659,
    20.73227, 25.04635, 29.9826, 35.39877, 41.64613, 49.05471, 55.54793,
    60.2282, 63.80492, 65.71034, 66.27112, 66.28201, 66.10315, 66.89112,
    66.59531, 64.6897,
  6.389893, 5.478107, 6.064652, 6.22161, 6.351696, 6.325079, 6.50585,
    6.656675, 6.769559, 7.338526, 8.694227, 10.86769, 14.07811, 17.54309,
    21.48107, 26.16568, 31.76213, 37.48363, 43.79842, 50.68221, 56.51512,
    60.86951, 64.28825, 65.76989, 66.0835, 65.79758, 65.31534, 65.90202,
    65.90208, 63.90043,
  6.410616, 5.452073, 6.06368, 6.240873, 6.511833, 6.751698, 7.09848,
    7.484078, 7.855348, 8.389054, 9.440147, 10.84754, 12.72334, 16.1798,
    20.35304, 25.16213, 30.55503, 36.98005, 43.39857, 50.76162, 56.87946,
    61.58752, 64.64639, 66.1299, 66.19158, 65.51664, 65.37741, 65.51433,
    64.89493, 60.73767,
  7.113036, 5.865105, 6.403191, 6.460069, 6.620265, 7.014742, 7.341809,
    6.453064, 6.338483, 7.339964, 8.757721, 10.76928, 13.33496, 16.58233,
    20.61019, 25.03129, 30.57186, 37.02738, 43.93519, 50.88341, 57.22113,
    62.00216, 65.00156, 66.22835, 66.05225, 65.79639, 65.96631, 65.55972,
    64.25658, 61.07912,
  9.64365, 7.746094, 7.72217, 7.472452, 7.319553, 7.191349, 6.260279,
    6.211018, 6.610363, 7.537637, 9.181958, 11.42267, 14.00761, 17.38088,
    21.35473, 25.11943, 30.40465, 37.43351, 44.77311, 51.65414, 57.84073,
    62.58061, 65.23088, 65.98542, 65.82565, 66.16852, 66.08925, 65.08157,
    61.17976, 61.64009,
  14.05975, 11.90847, 10.81475, 9.839365, 9.44438, 8.553796, 6.745733,
    7.010614, 7.081512, 7.843793, 9.549878, 12.51084, 15.50524, 18.0602,
    21.1787, 25.68591, 31.04846, 37.28317, 44.23098, 51.69415, 58.40272,
    62.94423, 64.7092, 64.89243, 65.29836, 65.74041, 65.43729, 63.87353,
    60.91351, 60.64587,
  18.4327, 15.63886, 15.79378, 13.69757, 12.70045, 11.11867, 9.628686,
    8.752954, 8.637225, 9.489635, 10.79951, 13.20156, 15.4119, 18.56609,
    22.39466, 26.46199, 31.44166, 37.23781, 43.7203, 50.7148, 58.07066,
    62.72072, 64.43244, 64.79739, 65.29369, 65.01904, 63.88723, 61.45367,
    61.89558, 60.76822,
  18.89345, 16.30091, 18.96247, 19.26081, 18.22838, 14.95948, 12.09188,
    9.526449, 8.62534, 9.351274, 10.93275, 13.22631, 16.55163, 19.35684,
    22.73621, 27.61959, 32.16249, 37.96112, 44.35616, 50.8211, 57.22224,
    62.47525, 64.26263, 65.19852, 65.51633, 64.6878, 61.57013, 63.63428,
    62.6372, 61.48045,
  10.00965, 10.80734, 12.96266, 15.75493, 17.83837, 17.55202, 12.01042,
    7.482879, 10.97987, 10.20076, 11.99634, 13.57981, 16.19187, 19.21564,
    22.96386, 26.84963, 32.29681, 38.3581, 44.88104, 51.61403, 57.6255,
    61.95395, 64.13596, 64.32327, 64.33257, 64.01723, 62.4444, 63.47438,
    63.36532, 62.39199,
  6.744746, 5.238547, 5.440132, 5.633987, 6.19508, 6.964653, 7.934439,
    9.162787, 8.562354, 9.937966, 12.13419, 14.75139, 17.09303, 19.6096,
    23.45526, 27.45336, 31.66, 38.62919, 45.67772, 52.32256, 57.49198,
    61.49556, 63.33836, 63.77089, 62.01286, 62.20988, 61.76054, 61.42893,
    61.67358, 61.72163,
  7.561798, 6.259003, 6.842371, 6.869125, 7.119063, 7.200011, 7.486839,
    7.768025, 8.451321, 10.18049, 12.4114, 15.07, 17.75225, 20.79307,
    23.55385, 26.95305, 32.41111, 37.02335, 44.55973, 51.91423, 56.89701,
    60.83603, 62.61618, 63.04612, 63.43273, 62.63098, 61.97107, 61.50953,
    61.07355, 60.93935,
  6.474945, 5.646083, 6.243909, 6.460885, 6.879009, 7.380854, 8.019196,
    8.485114, 9.257786, 11.37988, 14.38916, 17.00117, 19.63783, 21.60327,
    24.54758, 28.2519, 32.07213, 37.00153, 44.32853, 51.4964, 56.47479,
    60.73612, 62.3907, 63.17463, 63.31684, 62.70847, 61.91124, 61.47193,
    61.04987, 60.91547,
  6.130392, 4.735907, 5.326192, 5.519363, 5.92154, 6.369209, 6.909045,
    7.669654, 9.043941, 11.34749, 14.20438, 17.47927, 21.37238, 24.05401,
    27.0634, 30.23667, 33.8818, 38.97133, 46.22578, 52.40237, 57.08478,
    61.0336, 62.74501, 63.26826, 63.29988, 62.86217, 61.91653, 61.03177,
    60.77333, 60.82264,
  8.613836, 5.964026, 5.455208, 5.166882, 5.535852, 5.690979, 6.039802,
    6.535151, 7.45921, 9.046443, 12.02301, 15.80187, 19.63688, 24.88611,
    29.16553, 32.51451, 36.32311, 42.0565, 49.11222, 55.21351, 58.62653,
    61.8642, 63.36125, 63.88209, 63.17137, 62.59042, 61.93123, 60.88653,
    60.62605, 60.69139,
  16.81221, 11.49636, 7.6565, 4.098503, 5.518476, 5.346321, 5.64082,
    6.062425, 6.835322, 8.212239, 10.48968, 13.38156, 16.87106, 21.63329,
    27.52716, 32.47106, 37.91916, 45.02034, 53.08973, 59.34747, 62.63594,
    63.92384, 64.50691, 65.02798, 63.93361, 63.07014, 62.25463, 61.04301,
    60.58498, 60.72522,
  16.68628, 11.80449, 7.76299, 4.620072, 5.67802, 5.561226, 5.845536,
    6.277859, 7.231894, 8.827732, 10.82673, 12.77454, 15.8778, 19.93047,
    24.58302, 29.76189, 35.91096, 43.02795, 51.04397, 57.71265, 62.50981,
    64.82819, 65.26437, 65.49451, 65.03281, 63.50402, 62.4943, 61.24878,
    60.56465, 60.73115,
  17.45255, 12.80787, 8.736243, 5.958111, 6.688634, 6.55369, 6.796593,
    7.165847, 8.080982, 9.605744, 11.48289, 13.71078, 16.81728, 20.23008,
    24.64563, 29.7057, 35.70285, 42.67014, 49.91796, 56.38737, 61.30077,
    64.54374, 65.77302, 65.66388, 65.09082, 63.96025, 62.46583, 61.23387,
    60.56895, 60.73211,
  18.25648, 14.2444, 10.16702, 7.826877, 8.823427, 8.77292, 9.115061,
    9.441784, 10.33557, 11.63607, 13.21471, 15.70388, 19.00854, 22.53652,
    26.67007, 31.59572, 37.40682, 43.92945, 50.33695, 56.30985, 61.25524,
    64.40793, 65.8846, 65.99354, 65.41573, 64.51596, 62.77649, 61.64905,
    60.67813, 60.7389,
  18.5381, 15.03519, 11.43468, 9.398643, 10.83581, 11.37568, 12.04882,
    12.62735, 13.69304, 15.00977, 16.83798, 19.71125, 23.09442, 26.74939,
    30.6769, 35.44417, 41.10092, 47.08114, 53.07691, 58.16567, 62.45131,
    65.12344, 66.14707, 66.25626, 66.0472, 65.08537, 63.94322, 62.46486,
    61.372, 60.83397,
  18.54735, 15.00439, 11.87995, 10.12643, 11.37607, 11.99966, 13.21369,
    14.69537, 16.54471, 18.0629, 20.31616, 24.16047, 28.56847, 32.56467,
    36.03717, 40.43246, 45.6015, 51.28171, 56.83604, 61.82811, 65.54368,
    67.38744, 67.52423, 67.16685, 66.9409, 66.29078, 65.14969, 63.69206,
    62.45779, 61.52883,
  18.15535, 13.88316, 10.69942, 8.583516, 9.771317, 10.42335, 11.75561,
    13.62569, 15.69368, 17.30618, 19.61045, 23.65693, 28.4259, 32.61332,
    36.03066, 40.491, 45.58308, 51.29171, 57.15847, 62.57349, 66.52652,
    68.38618, 68.19026, 67.34605, 67.23496, 66.74117, 65.85055, 64.28271,
    63.1612, 62.32911,
  20.4035, 16.29085, 12.87685, 10.76204, 11.58429, 12.11468, 13.61763,
    15.70417, 17.41146, 18.93735, 21.70603, 25.5038, 30.01603, 33.80261,
    36.95073, 41.1446, 45.89608, 51.09858, 56.69331, 62.25477, 66.45277,
    68.59195, 68.54219, 67.91927, 67.61271, 66.8177, 66.0164, 64.56654,
    62.77433, 61.80937,
  30.48425, 26.828, 23.48429, 21.35666, 22.23756, 22.52691, 23.86055,
    25.42164, 26.73221, 28.24965, 30.79964, 34.09481, 37.98493, 41.06712,
    43.44764, 46.58348, 50.07717, 54.1318, 58.56295, 63.07761, 66.63891,
    68.58529, 68.85639, 68.3588, 68.02895, 67.27432, 66.58518, 65.29993,
    63.60765, 61.46349,
  46.1562, 44.39439, 41.7353, 40.42397, 41.36617, 41.78097, 42.58774,
    43.37585, 43.88247, 44.64082, 45.82925, 47.74751, 50.29031, 52.36656,
    53.65097, 55.29856, 56.99589, 59.09507, 61.81705, 64.73251, 66.78313,
    67.74713, 67.68144, 67.25853, 67.19804, 66.73125, 66.04946, 65.27238,
    64.46376, 62.90473,
  54.85276, 55.22938, 55.51852, 56.26041, 57.10941, 58.11211, 58.33539,
    58.16706, 58.1197, 58.1375, 58.07431, 58.0481, 58.24078, 58.8605,
    59.31526, 59.92151, 60.62005, 61.49524, 62.40101, 63.36356, 64.54356,
    65.66293, 66.106, 65.80843, 65.73813, 65.44169, 64.92427, 64.15063,
    63.80181, 62.91941,
  62.6137, 62.60626, 62.60863, 62.69595, 63.27102, 64.23483, 64.79514,
    64.40257, 63.79419, 63.98265, 64.01671, 63.9366, 63.59776, 63.30451,
    63.15361, 63.1227, 63.07409, 62.29295, 62.22507, 62.33022, 62.05419,
    62.82757, 63.61922, 63.95034, 63.97196, 64.2579, 63.97727, 62.82236,
    61.71583, 60.94326,
  20.68032, 23.33181, 26.10992, 28.9422, 32.20782, 35.57121, 39.00137,
    42.58931, 46.38411, 49.96664, 53.81118, 57.2224, 59.86152, 61.8475,
    63.1272, 63.76419, 63.91963, 63.82161, 63.48501, 62.83347, 61.6843,
    60.05638, 58.36951, 56.83346, 55.33391, 53.93757, 53.26947, 53.64528,
    52.96299, 51.74152,
  19.49576, 22.27382, 25.64359, 28.79585, 32.26164, 36.01258, 39.80918,
    43.70994, 47.53531, 51.21909, 54.98169, 58.56124, 61.47795, 63.34179,
    64.20387, 64.52457, 64.47249, 64.28254, 63.99217, 63.5899, 62.76379,
    61.52812, 59.90916, 58.3568, 57.01836, 55.27891, 53.52942, 53.29727,
    52.82339, 51.95933,
  20.10416, 22.60864, 25.83496, 29.217, 32.50402, 36.13968, 40.00023,
    44.15708, 48.33543, 52.15335, 55.66287, 59.02664, 61.87157, 63.8703,
    64.85338, 64.90169, 64.56071, 64.1795, 63.7349, 63.19322, 62.7336,
    61.83133, 60.35821, 58.68132, 57.19715, 56.29125, 55.54978, 53.88017,
    52.75783, 51.49539,
  21.18771, 23.67125, 27.26155, 30.13522, 33.37519, 36.55714, 40.09332,
    44.18893, 48.52545, 52.72926, 56.35794, 59.59027, 62.43888, 64.33898,
    65.39955, 65.69501, 65.1487, 64.39016, 63.95069, 63.42475, 62.79457,
    61.36053, 59.12518, 57.83941, 56.40461, 56.23539, 56.4436, 55.79428,
    54.0468, 52.88622,
  22.11494, 24.91681, 28.16483, 31.71662, 34.58957, 37.48782, 40.40885,
    44.25093, 48.11244, 52.37896, 56.30173, 59.7133, 62.80962, 64.94965,
    66.11134, 66.40157, 65.84219, 64.92228, 64.29512, 63.58959, 62.35509,
    60.46164, 58.79622, 57.43974, 56.18514, 55.53093, 55.48641, 56.62712,
    56.34995, 53.90481,
  23.17372, 25.48859, 28.93611, 32.393, 35.87035, 38.77116, 41.36665,
    45.31568, 48.75552, 52.09909, 55.7848, 59.39161, 62.76184, 64.96975,
    66.40379, 66.95381, 66.2951, 65.52538, 64.40733, 63.50351, 62.10192,
    59.97989, 58.96844, 57.58515, 56.32895, 55.4348, 54.84624, 55.48402,
    55.52923, 52.77266,
  26.06911, 27.3373, 29.83167, 32.86994, 36.25131, 39.45148, 42.48013,
    46.25531, 50.01569, 53.24091, 56.50353, 59.08595, 60.77132, 63.02403,
    64.356, 65.14775, 65.31266, 64.58479, 63.29735, 62.42198, 61.26655,
    59.89659, 58.66063, 57.60792, 56.39609, 55.42046, 55.21619, 55.20362,
    54.36074, 50.14907,
  31.03424, 31.54531, 32.87373, 34.74313, 37.42189, 40.75568, 43.95578,
    45.95021, 48.76994, 52.16278, 55.24897, 57.99686, 60.57038, 62.70734,
    64.1254, 64.77109, 65.20982, 65.09063, 64.13502, 62.74134, 61.26801,
    59.74255, 58.33969, 57.14256, 56.03202, 55.51666, 55.60236, 55.02953,
    53.33573, 50.46709,
  36.43989, 37.76844, 38.22355, 38.98812, 40.1848, 42.44466, 43.89463,
    46.66745, 50.13866, 53.29328, 56.11086, 58.49984, 60.48626, 62.3681,
    63.83877, 64.22802, 64.69685, 65.24691, 65.19315, 63.85794, 61.99795,
    60.02058, 58.18602, 56.43403, 55.35299, 55.44193, 55.41179, 54.27911,
    50.30777, 51.00761,
  39.17206, 42.71449, 44.49768, 45.04723, 45.00146, 45.33929, 45.65199,
    48.04019, 50.93431, 54.209, 56.83667, 59.13158, 60.65592, 61.7999,
    62.48215, 63.26741, 63.68753, 64.02065, 64.10725, 63.53049, 62.6225,
    60.39546, 57.95906, 55.84425, 54.98998, 54.71066, 54.28905, 52.7279,
    50.58234, 50.21584,
  37.88478, 41.26136, 46.33141, 49.18928, 50.18029, 49.81503, 49.89831,
    50.8084, 52.33744, 55.59529, 57.72991, 59.12793, 60.39288, 61.44624,
    62.14843, 62.54975, 62.66673, 62.62151, 62.51479, 62.17707, 62.11078,
    60.41993, 57.70041, 56.10938, 55.50403, 54.43232, 52.74597, 51.83913,
    51.65119, 50.52347,
  34.69719, 35.03256, 42.43894, 48.58686, 54.22822, 54.17727, 52.57893,
    51.74854, 53.84888, 55.90745, 58.42339, 59.96862, 61.73238, 62.62573,
    62.93042, 62.90409, 63.04432, 62.87886, 62.30542, 61.44605, 61.18075,
    60.17551, 57.49466, 55.89172, 55.18075, 54.05787, 50.59541, 52.50978,
    52.3587, 51.37691,
  29.08014, 32.1901, 35.29385, 41.3245, 48.33426, 53.81057, 52.75154,
    50.63033, 56.73896, 57.85236, 60.39826, 61.91505, 63.39826, 64.4623,
    64.59077, 63.20556, 63.30569, 63.33757, 62.74197, 61.42469, 60.61861,
    59.43188, 57.44428, 55.22406, 53.76458, 53.01627, 51.51117, 52.24373,
    52.38947, 52.16625,
  27.14139, 29.78423, 32.30094, 35.43781, 39.03903, 42.92229, 48.06996,
    53.10754, 55.27215, 58.4932, 61.47565, 63.84906, 65.00079, 65.9495,
    65.92033, 64.58856, 63.6835, 63.54603, 63.403, 61.70302, 59.66109,
    58.05822, 56.07259, 54.63354, 52.16068, 51.49312, 51.48027, 50.66279,
    50.96255, 51.35402,
  25.55078, 27.34741, 31.2032, 35.23331, 38.86345, 42.95844, 46.3848,
    50.22523, 54.80659, 58.48177, 61.1738, 63.29033, 65.19836, 66.49831,
    66.62891, 66.56714, 65.01184, 63.71864, 62.84216, 61.60184, 58.95848,
    57.36165, 55.45183, 54.09515, 53.29818, 52.41416, 51.61819, 51.12936,
    50.51012, 50.35831,
  26.02097, 27.76018, 30.57687, 33.27625, 37.02176, 40.33297, 44.4239,
    48.27275, 52.52267, 57.03397, 60.45234, 62.91512, 65.05333, 66.8925,
    67.47743, 67.1219, 66.76331, 65.23815, 63.63685, 61.83316, 59.80925,
    57.96907, 55.58128, 54.01006, 53.22599, 52.41864, 51.32946, 50.87956,
    50.57174, 50.445,
  27.89702, 28.68701, 31.63808, 34.4417, 37.62928, 40.81825, 44.16247,
    47.24144, 50.84476, 55.05939, 58.76213, 61.93139, 64.83672, 66.45464,
    67.48846, 68.07484, 68.35744, 67.87318, 66.04508, 63.47831, 60.55313,
    58.70787, 56.49676, 54.53603, 53.32904, 52.66857, 51.39222, 50.50806,
    50.32825, 50.34461,
  34.65483, 32.95899, 33.70572, 35.7668, 39.49212, 42.72883, 45.79095,
    49.0746, 51.83281, 55.1073, 58.52786, 61.64518, 63.53453, 64.99733,
    65.97106, 67.14271, 68.53872, 69.34277, 68.90022, 66.66819, 62.94945,
    59.67044, 57.40957, 55.58838, 53.85503, 52.75994, 51.67941, 50.43645,
    50.21812, 50.24089,
  44.87836, 41.83962, 38.29705, 36.79692, 41.17216, 44.22746, 47.88735,
    50.95203, 54.57405, 57.57076, 60.46975, 62.5373, 63.85796, 64.50977,
    64.61145, 65.32747, 66.69044, 68.05964, 68.36289, 67.81868, 65.52831,
    61.46194, 58.15461, 56.57147, 54.6137, 53.71646, 52.40022, 50.71273,
    50.17316, 50.25442,
  44.8251, 42.99033, 39.67625, 38.48711, 42.63192, 45.66071, 49.49177,
    53.12881, 56.67606, 59.94927, 62.66786, 64.35688, 65.91235, 66.57765,
    66.5067, 65.99419, 65.95911, 66.11697, 65.56161, 64.8901, 64.06837,
    62.02842, 58.89311, 56.7086, 55.0973, 54.00902, 52.86901, 51.01017,
    50.14899, 50.28191,
  46.68955, 44.578, 41.48388, 40.564, 44.64957, 47.59997, 51.46059, 55.35725,
    59.09179, 62.52606, 64.98331, 66.65501, 68.21651, 68.99934, 68.99673,
    68.63797, 67.98437, 67.16824, 66.00095, 64.22131, 62.88088, 61.53148,
    59.43608, 56.94732, 55.21663, 54.01808, 52.86329, 51.25335, 50.17543,
    50.28574,
  50.75454, 48.75051, 45.35391, 44.31499, 48.54078, 51.27822, 54.8292,
    58.36737, 62.1836, 65.80328, 68.58083, 70.53315, 71.83035, 72.28444,
    72.07351, 71.39021, 70.27966, 69.01319, 67.43118, 65.52462, 63.63697,
    61.8055, 59.93027, 57.44088, 55.61604, 54.03828, 53.06664, 51.86985,
    50.59404, 50.29081,
  58.47437, 56.04452, 52.55104, 50.93638, 54.45876, 57.10823, 60.25652,
    63.349, 66.52567, 69.65627, 72.72546, 75.49208, 77.36571, 77.76582,
    77.09422, 76.18459, 74.70094, 72.78888, 70.54295, 68.2204, 66.08488,
    63.38002, 60.73174, 58.07808, 56.47369, 54.76824, 53.37836, 52.52332,
    51.62159, 50.59473,
  68.06389, 65.15018, 61.40654, 59.19145, 61.35235, 62.68797, 65.2342,
    68.00769, 71.16792, 73.4922, 75.8578, 79.06567, 82.22272, 83.32523,
    82.27431, 81.32265, 79.81789, 77.7591, 74.93321, 72.38374, 69.8465,
    66.41349, 62.36438, 59.3927, 57.7784, 56.23657, 54.55598, 52.87534,
    52.30048, 51.49813,
  74.83125, 71.27983, 66.21134, 63.37344, 64.49356, 64.81857, 66.34337,
    68.65561, 71.39627, 72.84392, 74.33991, 76.94308, 79.95834, 81.14858,
    80.14859, 79.71133, 78.64188, 77.27454, 75.05057, 72.72182, 70.49036,
    67.27251, 63.01718, 59.80307, 58.25027, 56.92284, 55.44919, 53.3776,
    52.30964, 52.04974,
  75.61665, 71.36346, 66.35155, 63.03781, 63.48376, 63.25626, 64.3847,
    66.17608, 67.77837, 68.21626, 69.8106, 72.12976, 75.08767, 76.18387,
    75.10882, 74.74837, 74.10143, 72.97474, 71.60381, 70.20253, 68.43994,
    66.13758, 62.51525, 59.75035, 58.37346, 56.88829, 55.66562, 53.89481,
    52.30877, 51.51375,
  70.76257, 67.38416, 62.82854, 59.84638, 60.33044, 59.81321, 60.31363,
    61.34802, 61.86816, 61.74462, 62.66319, 64.61814, 67.46127, 68.94389,
    68.41964, 68.21422, 67.6868, 67.10861, 66.02233, 65.33727, 64.38729,
    63.11779, 60.87666, 58.89814, 58.05352, 56.72569, 55.76762, 54.36048,
    52.84837, 51.54024,
  62.61716, 60.68987, 57.9538, 56.16518, 56.73803, 56.77968, 57.00924,
    57.49239, 57.45194, 57.06828, 56.85823, 57.61188, 59.3695, 60.72353,
    60.72603, 60.69081, 60.65586, 60.29902, 59.92569, 59.96202, 59.90949,
    59.32187, 57.98359, 56.88465, 56.60445, 55.94867, 54.95936, 53.9062,
    53.25795, 52.68618,
  53.01891, 53.0147, 53.06205, 53.3949, 53.74717, 54.28151, 54.46734,
    54.56975, 54.68233, 54.53323, 54.20641, 53.67693, 53.30621, 53.63096,
    53.70984, 53.71819, 53.79504, 53.91998, 53.92569, 53.95124, 54.33738,
    55.01486, 55.29436, 54.94131, 54.95115, 54.59538, 53.9418, 53.07162,
    52.55819, 52.12275,
  52.93715, 52.73519, 52.59219, 52.51409, 52.79576, 53.27539, 53.64447,
    53.57507, 53.12456, 53.63281, 53.6686, 53.46194, 52.99378, 52.72446,
    52.65619, 52.62158, 52.49884, 51.72018, 51.28759, 51.28836, 51.04645,
    51.65166, 52.54866, 52.99583, 53.02284, 53.29627, 53.18961, 52.22383,
    51.01608, 50.39513,
  55.20652, 57.04173, 57.92033, 58.75338, 59.21657, 59.50416, 59.47416,
    59.21326, 58.64933, 57.94523, 57.27731, 56.68038, 55.99259, 55.35358,
    54.81172, 54.37935, 54.12668, 53.95844, 53.92204, 53.82504, 53.35313,
    52.60997, 51.86768, 51.33071, 50.82349, 50.06613, 49.6793, 49.88182,
    49.49212, 47.99209,
  55.37307, 57.16596, 58.07474, 59.02233, 59.53763, 59.75012, 59.69005,
    59.62193, 59.18416, 58.55593, 57.75008, 57.04045, 56.44904, 55.71285,
    54.96118, 54.45918, 54.10016, 53.97157, 54.02251, 54.06596, 54.03684,
    53.74911, 53.3061, 52.91887, 52.36817, 51.02863, 49.64251, 49.47778,
    49.17945, 48.0643,
  55.43731, 57.13029, 57.9118, 58.87671, 59.48773, 59.71836, 59.6081,
    59.44007, 59.16901, 58.62121, 58.00263, 57.35945, 56.6393, 55.90781,
    55.25819, 54.54068, 54.02047, 53.79094, 53.65462, 53.66489, 53.79605,
    53.96567, 53.89183, 53.46682, 52.98383, 52.1718, 51.27181, 49.94332,
    49.1697, 47.91054,
  55.69445, 57.18188, 57.88288, 58.8606, 59.55667, 59.94532, 59.92389,
    59.67546, 59.20428, 58.57753, 58.08293, 57.92512, 57.35394, 56.36153,
    55.624, 55.0983, 54.53234, 53.98135, 53.76896, 53.71146, 53.71554,
    53.38044, 52.46573, 52.64016, 52.29793, 52.57458, 52.49714, 51.7568,
    50.57102, 49.76857,
  55.90132, 57.33447, 57.93614, 58.69482, 59.25737, 59.74001, 60.08955,
    59.89372, 59.36673, 58.47945, 58.00739, 58.22346, 58.24729, 57.32076,
    56.36037, 55.68366, 55.07962, 54.54058, 54.25879, 53.93306, 53.3425,
    52.6019, 52.05437, 52.06951, 52.11322, 51.94907, 52.12057, 53.02889,
    52.8192, 50.85661,
  56.51961, 57.71415, 58.37392, 58.90965, 59.09996, 59.46056, 60.06084,
    60.23817, 59.8641, 59.14737, 58.67808, 58.6484, 58.70876, 57.85979,
    57.12823, 56.3689, 55.32458, 54.86455, 54.52438, 54.228, 53.42041,
    52.24067, 52.32399, 52.15616, 51.98191, 51.78488, 51.48227, 52.03074,
    52.04319, 49.74327,
  58.35777, 58.71692, 59.25002, 59.47063, 59.495, 59.67342, 60.101, 60.04517,
    59.77936, 59.13285, 58.7795, 57.97538, 56.66663, 56.26762, 55.60716,
    55.13995, 54.80223, 54.0059, 53.25894, 52.96268, 52.54908, 52.21665,
    52.16594, 52.24449, 52.0263, 51.82989, 51.84019, 51.84382, 51.04606,
    46.89738,
  62.34925, 61.42764, 60.94668, 60.64913, 60.37293, 60.50333, 60.4319,
    58.99717, 57.70933, 57.29097, 56.84366, 56.4996, 56.28094, 55.95919,
    55.63854, 55.35033, 55.05696, 54.5793, 53.90022, 53.20322, 52.52486,
    52.10144, 51.92126, 51.89917, 51.84197, 52.00215, 52.16184, 51.48083,
    50.22417, 47.13623,
  67.4622, 66.70174, 64.60315, 63.13255, 62.12342, 61.30375, 59.64255,
    59.22333, 58.46625, 57.47332, 56.79331, 56.29757, 55.6952, 55.36995,
    55.19686, 54.83834, 54.92296, 55.11826, 54.99167, 54.16043, 53.2665,
    52.41896, 51.76382, 51.25619, 51.17645, 51.86444, 52.08037, 50.99451,
    47.04573, 47.60288,
  70.1036, 71.90245, 70.40459, 68.21906, 65.87103, 63.31808, 60.42937,
    60.02646, 59.22424, 58.29303, 56.91351, 55.96686, 55.11572, 54.34653,
    53.84831, 53.85129, 53.91141, 54.17506, 54.37741, 54.1414, 53.86182,
    52.81312, 51.73155, 50.93196, 50.99139, 51.15319, 50.97934, 49.65348,
    47.19356, 47.16465,
  67.84053, 70.80186, 74.03661, 73.59724, 71.59726, 67.15922, 63.7085,
    61.43363, 59.95173, 59.55437, 57.64587, 55.68446, 54.79722, 54.04483,
    53.39666, 53.11202, 52.95104, 52.91404, 53.11008, 53.20302, 53.40385,
    52.6611, 51.51172, 51.26771, 51.65252, 51.24129, 49.7168, 48.1037,
    48.24269, 47.34156,
  63.85205, 64.38001, 69.47006, 73.52002, 74.45542, 71.27387, 66.71778,
    62.75093, 61.00985, 60.05426, 58.5636, 57.13431, 56.18005, 55.37069,
    54.23536, 53.44478, 53.32852, 53.1473, 52.91144, 52.66664, 52.87034,
    52.41035, 51.21677, 50.86693, 51.16475, 50.76275, 47.48413, 49.56673,
    49.15064, 48.00853,
  58.49988, 60.47489, 61.83953, 64.86962, 67.96079, 69.54698, 65.37749,
    61.64375, 63.43931, 61.76329, 60.56286, 58.89235, 58.04825, 57.13969,
    55.70691, 53.7366, 53.67477, 53.68535, 53.42715, 52.80142, 52.67755,
    52.23387, 51.21049, 50.18122, 49.77578, 49.78431, 47.87201, 49.30066,
    49.43584, 48.70559,
  59.21059, 60.12395, 59.9602, 59.03988, 58.66085, 59.90353, 61.80134,
    62.87255, 61.14047, 61.78791, 61.56209, 60.19897, 59.10831, 58.18053,
    56.51563, 54.77395, 53.88893, 53.89211, 54.02863, 53.15284, 52.28786,
    51.41078, 50.25087, 49.6529, 47.54786, 47.77109, 48.05597, 47.42123,
    47.60755, 47.97107,
  59.63934, 60.74486, 61.20815, 61.25539, 61.02663, 60.75977, 60.89425,
    60.64095, 60.1023, 59.63412, 59.46273, 59.00575, 58.80478, 58.21212,
    57.05753, 56.23025, 54.7328, 53.87109, 53.48956, 52.79601, 51.33761,
    50.68536, 49.76232, 48.88524, 49.36919, 48.60556, 48.14846, 47.68822,
    47.24692, 47.15115,
  60.11044, 61.25177, 61.71618, 61.82301, 61.53123, 61.52647, 61.51297,
    61.18695, 60.12845, 59.05829, 58.60598, 58.55171, 58.67648, 59.05,
    58.14159, 56.85433, 56.18438, 55.02164, 53.89035, 52.84241, 51.74141,
    50.84681, 49.77618, 49.38796, 49.13245, 48.59934, 47.94477, 47.5541,
    47.31514, 47.25545,
  62.68132, 62.94823, 63.28059, 63.50487, 63.10769, 62.34498, 61.91597,
    61.99059, 61.30358, 60.04025, 58.80819, 58.54174, 58.97274, 58.82475,
    58.54482, 58.30283, 57.99681, 57.41446, 56.05729, 54.29019, 52.43598,
    51.49687, 50.49459, 49.81385, 49.59393, 49.01017, 47.93183, 47.31884,
    47.17275, 47.19831,
  69.01507, 67.12213, 65.4722, 65.13634, 65.30071, 64.4823, 63.90569,
    63.17717, 62.8333, 61.52069, 60.44194, 59.47654, 58.45456, 57.50842,
    57.11821, 57.68539, 58.5139, 59.03571, 58.72877, 57.15042, 54.60622,
    52.46313, 51.44187, 50.77257, 50.06721, 49.25137, 48.24493, 47.20438,
    47.10477, 47.10789,
  78.50069, 74.51298, 69.28656, 66.08846, 67.4437, 66.76748, 65.957,
    65.14329, 63.97567, 63.09885, 62.19295, 61.0615, 59.34365, 57.5253,
    55.73655, 55.87107, 56.85334, 58.06713, 58.65061, 58.58601, 56.98886,
    54.19659, 52.2602, 51.89963, 51.0377, 50.27863, 49.00383, 47.43048,
    47.10141, 47.15617,
  77.25568, 74.19534, 69.12437, 66.543, 68.00198, 68.03948, 67.71329,
    66.75856, 65.72504, 64.60902, 63.58677, 62.67289, 61.81127, 59.71587,
    57.7765, 56.44868, 56.19392, 56.52708, 56.39766, 56.20097, 55.76101,
    54.58635, 52.81285, 52.04396, 51.41324, 50.7975, 49.43718, 47.76777,
    47.06896, 47.18645,
  75.86208, 72.64543, 67.9217, 65.30566, 67.02025, 67.46013, 67.83704,
    67.65282, 67.29792, 66.40942, 65.1664, 63.81599, 62.95744, 61.85435,
    60.15947, 58.97096, 58.21426, 57.6945, 57.01222, 55.86172, 54.95743,
    54.35894, 53.51141, 52.23391, 51.48418, 50.71293, 49.57817, 48.01425,
    47.02956, 47.12279,
  73.25181, 70.70763, 65.38392, 63.06408, 64.73933, 65.37164, 66.41902,
    67.05627, 67.84283, 68.27106, 67.42746, 66.08543, 65.0017, 63.90125,
    62.54767, 61.24999, 60.19891, 59.33935, 58.33714, 57.04961, 55.71864,
    54.69426, 54.17046, 52.6707, 51.75317, 50.80548, 50.08104, 48.65034,
    47.35366, 47.11991,
  70.60606, 68.09056, 63.28357, 60.80869, 62.38807, 63.09567, 64.46904,
    65.64222, 67.27367, 68.54932, 69.1161, 68.98215, 68.81295, 68.21657,
    66.87528, 65.65517, 64.25298, 62.83517, 61.26644, 59.65255, 58.06608,
    56.28479, 55.14679, 53.56263, 52.67905, 51.61082, 50.44646, 49.50558,
    48.25621, 47.37616,
  68.50005, 65.19768, 61.42585, 58.88065, 60.08318, 60.5621, 62.09525,
    64.09994, 66.2784, 67.81633, 68.95564, 70.77059, 72.67834, 73.11285,
    71.88411, 70.86593, 69.26901, 67.49873, 65.4226, 63.57805, 61.72998,
    59.51218, 56.83724, 55.15133, 54.32618, 53.15672, 51.54017, 49.88781,
    49.04743, 48.10616,
  67.28165, 63.72716, 58.7578, 56.48858, 57.07336, 57.39806, 59.04692,
    61.44936, 64.04999, 64.74303, 65.73273, 67.92862, 70.53181, 71.56137,
    70.47747, 69.8732, 68.97489, 67.67687, 66.00186, 64.40282, 62.53168,
    60.28724, 57.42281, 55.44703, 54.76035, 53.62246, 52.35548, 50.31547,
    49.19979, 48.48532,
  66.38506, 62.55197, 58.19064, 55.19408, 55.61573, 55.43242, 56.6199,
    58.80769, 60.68488, 60.95093, 62.38605, 64.75911, 67.50687, 68.50127,
    67.49894, 67.10221, 66.57393, 65.63684, 64.46605, 63.51451, 62.05069,
    60.04013, 57.39154, 55.42159, 54.79644, 53.55901, 52.38148, 50.80539,
    49.30545, 48.17239,
  63.61885, 60.73564, 56.75305, 54.20348, 54.62144, 54.18829, 54.7836,
    55.91879, 56.82053, 56.85284, 57.79427, 59.89405, 62.62321, 63.98074,
    63.19467, 62.97583, 62.81079, 62.28109, 61.37312, 60.82062, 60.03125,
    58.78774, 56.70699, 55.23455, 54.71941, 53.64833, 52.61027, 51.12758,
    49.77241, 48.15152,
  58.38933, 56.79167, 54.13574, 52.34591, 52.97454, 53.01719, 53.15709,
    53.69692, 53.87913, 53.5035, 53.43262, 54.40655, 56.21444, 57.57107,
    57.39851, 57.24301, 57.19279, 57.08632, 56.75732, 56.68454, 56.59384,
    55.98503, 54.61029, 53.66388, 53.58737, 52.95987, 52.01131, 50.92053,
    50.18029, 49.07714,
  49.80633, 49.89758, 49.9279, 50.16767, 50.54329, 51.09441, 51.36971,
    51.43303, 51.53388, 51.37425, 51.0322, 50.49028, 50.22081, 50.52803,
    50.65936, 50.72091, 50.75232, 50.86612, 50.89754, 51.01502, 51.37137,
    51.95541, 52.30472, 51.92281, 51.88411, 51.55003, 50.96727, 50.1867,
    49.32717, 48.7331,
  49.80103, 49.64721, 49.52517, 49.44127, 49.75069, 50.24334, 50.60138,
    50.62336, 49.98967, 50.19931, 50.44159, 50.35287, 49.86214, 49.62614,
    49.53785, 49.53253, 49.37266, 48.26216, 48.03805, 47.96325, 47.86565,
    48.50657, 49.51579, 50.00975, 49.92443, 50.05565, 49.75097, 48.80341,
    47.85794, 47.27098,
  53.81927, 53.39288, 53.14958, 52.93203, 52.63325, 52.40189, 52.18358,
    51.91237, 51.67396, 51.52534, 51.48307, 51.4363, 51.3, 51.28373,
    51.28748, 51.34021, 51.40561, 51.44481, 51.38366, 51.27997, 51.03497,
    50.64988, 50.41504, 50.34173, 50.20626, 49.6876, 46.73523, 48.41066,
    45.73882, 44.16094,
  54.23049, 53.84269, 53.47748, 53.21, 52.93021, 52.68996, 52.53385,
    52.30596, 52.03848, 51.81903, 51.65449, 51.59956, 51.55526, 51.36934,
    51.25368, 51.23395, 51.3037, 51.54626, 51.79472, 52.02914, 52.14065,
    52.10498, 51.91094, 51.78806, 51.40929, 50.08466, 48.05383, 46.388,
    45.36255, 44.2608,
  54.17259, 53.95513, 53.68136, 53.39998, 53.07175, 52.78414, 52.59713,
    52.44142, 52.24928, 52.02127, 51.92722, 51.90346, 51.80909, 51.72817,
    51.55962, 51.19032, 50.99967, 51.11456, 51.34357, 51.75756, 52.3889,
    52.92873, 53.04126, 52.80799, 52.13709, 51.103, 50.33568, 49.21451,
    44.84867, 44.26651,
  54.00097, 53.8115, 53.6722, 53.54364, 53.37436, 53.175, 52.89146, 52.66815,
    52.44146, 52.14651, 52.08627, 52.3475, 52.45227, 52.22286, 52.04564,
    51.80631, 51.4818, 51.22788, 51.25014, 51.50072, 52.07736, 52.23081,
    51.84406, 51.98554, 51.67437, 51.91113, 51.42215, 50.82364, 49.94925,
    46.01038,
  53.8784, 53.48431, 53.30993, 53.25845, 53.20968, 53.26188, 53.32282,
    53.02963, 52.65081, 52.1997, 52.19619, 52.7916, 53.24259, 52.96788,
    52.7028, 52.50946, 52.17162, 51.87056, 51.77409, 51.60984, 51.47958,
    51.40132, 51.2151, 51.50338, 51.51323, 51.26309, 51.34133, 52.18365,
    52.12623, 50.48529,
  54.08231, 53.59169, 53.20837, 52.91396, 52.79411, 53.08852, 53.6512,
    53.78996, 53.49435, 53.00062, 52.84043, 53.35974, 53.92369, 53.5519,
    53.31847, 53.04396, 52.28681, 52.13445, 52.23989, 52.11709, 51.69257,
    50.94376, 51.34573, 51.38074, 51.27128, 51.11533, 50.76608, 51.0566,
    51.22781, 49.61435,
  54.61287, 54.00252, 53.61319, 53.08091, 52.72077, 52.88976, 53.57431,
    53.88866, 53.99895, 53.63309, 53.49197, 53.04161, 52.07109, 52.10233,
    51.85326, 51.71734, 51.65416, 51.19955, 50.73519, 50.92801, 50.91327,
    50.93646, 51.27966, 51.61973, 51.58706, 51.42677, 51.40997, 51.24302,
    50.42934, 43.21169,
  56.07269, 54.77707, 54.29209, 53.72586, 53.237, 53.2468, 53.34716,
    52.30871, 51.6398, 51.72793, 51.81153, 51.87957, 52.05391, 52.17517,
    52.25377, 52.23597, 52.0274, 51.70041, 51.37368, 51.05156, 50.8287,
    50.78394, 51.00004, 51.35228, 51.4762, 51.74841, 51.80172, 51.12014,
    50.1158, 43.36165,
  59.50858, 57.47709, 55.85661, 54.87302, 54.18548, 53.55188, 52.21747,
    52.06649, 51.89297, 51.61656, 51.54469, 51.51486, 51.55553, 51.96,
    52.32484, 52.2471, 52.4586, 52.78186, 52.83658, 52.21673, 51.63201,
    51.11811, 50.86881, 50.58608, 50.77349, 51.63013, 51.93373, 50.71304,
    43.38467, 43.88767,
  63.7056, 62.58834, 60.07151, 57.95025, 56.64337, 54.74674, 52.5548,
    52.61315, 52.36359, 52.02061, 51.45874, 51.17757, 50.91017, 50.87373,
    50.90945, 51.31417, 51.7875, 52.31743, 52.5803, 52.56266, 52.42531,
    51.71889, 50.94233, 50.36621, 50.51271, 50.56995, 50.43363, 49.40795,
    43.37877, 43.4453,
  65.74505, 65.44868, 66.17703, 63.4956, 61.47732, 57.75169, 55.20038,
    53.65246, 52.89527, 52.98947, 51.82145, 50.71122, 50.43058, 50.27327,
    50.13546, 50.26095, 50.57776, 50.90461, 51.3465, 51.61225, 52.11753,
    51.68445, 50.86725, 50.9257, 51.55319, 51.12442, 49.46114, 43.97344,
    44.4928, 43.53173,
  64.31589, 63.58328, 66.62519, 68.1104, 66.51023, 62.62751, 58.48175,
    54.87523, 53.16293, 53.0384, 52.28776, 51.68159, 51.43765, 51.17453,
    50.64935, 50.36741, 50.57463, 50.81205, 51.00108, 51.14366, 51.6261,
    51.3604, 50.5739, 50.5206, 50.89922, 50.51934, 44.00705, 48.59557,
    45.20283, 44.1173,
  56.27878, 57.7434, 59.29353, 61.81131, 63.79266, 63.62035, 58.1128,
    53.65969, 55.65009, 54.04222, 53.49068, 52.75979, 52.6549, 52.4808,
    51.83416, 50.51238, 50.80628, 51.15678, 51.31669, 51.15925, 51.46071,
    51.37267, 50.66351, 49.87662, 49.59021, 49.47703, 44.26716, 46.12631,
    45.93365, 44.7257,
  55.71962, 54.81566, 54.30347, 53.1015, 52.87477, 53.80401, 55.10998,
    55.77826, 54.02966, 54.3139, 54.25783, 53.52026, 53.05774, 52.8667,
    52.10185, 51.1459, 50.88752, 51.42033, 51.8756, 51.35324, 50.93307,
    50.47072, 49.48779, 46.58605, 44.01373, 44.19486, 44.22726, 43.68088,
    43.96998, 44.12754,
  57.2611, 56.81971, 55.94675, 55.00208, 54.32479, 54.08462, 54.39107,
    54.42381, 53.91687, 53.55614, 53.2855, 52.87427, 52.84039, 52.55463,
    52.06195, 51.92426, 51.21679, 51.13369, 51.19755, 50.79528, 49.79109,
    49.51997, 48.01242, 44.60798, 45.51247, 45.00718, 44.46593, 43.88385,
    43.4328, 43.412,
  56.45895, 56.334, 55.91751, 55.23729, 54.66112, 54.55272, 54.57774,
    54.57777, 54.18259, 53.71386, 53.60738, 53.45213, 53.45045, 53.59544,
    52.73526, 51.97393, 51.85379, 51.45393, 51.02393, 50.41998, 49.30261,
    48.12339, 45.86859, 44.89693, 45.07874, 44.96183, 44.29548, 43.83015,
    43.5289, 43.51828,
  57.9109, 56.98038, 56.34727, 55.79876, 55.15762, 54.29121, 54.05784,
    54.35439, 54.25837, 53.94857, 53.76352, 54.22966, 54.96684, 54.81794,
    54.2306, 53.83687, 53.68225, 53.35917, 52.40926, 51.19596, 50.15659,
    49.11161, 46.8531, 45.43986, 45.4501, 45.26632, 44.28387, 43.59276,
    43.4503, 43.48758,
  62.53261, 59.8553, 57.7065, 56.73293, 56.25956, 55.41007, 54.91374,
    54.62288, 54.52714, 53.99192, 53.85195, 53.95965, 54.05716, 54.10154,
    54.24096, 54.80544, 55.46337, 55.83382, 55.39481, 53.87324, 51.98134,
    50.69075, 48.15654, 46.85981, 46.06548, 45.438, 44.43463, 43.48559,
    43.40377, 43.41094,
  71.81598, 66.86415, 61.06709, 57.49881, 57.89281, 56.98217, 56.43382,
    55.89863, 55.20272, 54.90424, 54.5597, 53.87172, 53.01861, 52.45832,
    52.03571, 52.72878, 54.08422, 55.65136, 56.44786, 56.20478, 54.67595,
    52.46094, 50.19466, 49.02971, 47.28039, 46.221, 45.06245, 43.73973,
    43.44381, 43.49302,
  71.12239, 67.41003, 61.95255, 58.97779, 59.43749, 58.88597, 58.38116,
    57.49178, 56.84425, 56.4873, 56.11666, 55.30247, 54.56479, 53.38364,
    52.29685, 51.73721, 52.063, 52.96267, 53.75368, 53.99695, 53.7704,
    52.90873, 51.8199, 50.34334, 48.58167, 46.75725, 45.52449, 44.07281,
    43.46665, 43.52008,
  70.78703, 67.69981, 62.39367, 59.96452, 60.82584, 60.64445, 60.40852,
    59.92297, 59.32387, 58.68927, 57.94475, 56.96094, 56.34256, 55.45323,
    54.40277, 53.70357, 53.38828, 53.44249, 53.44821, 52.95451, 52.5623,
    52.43119, 52.11611, 51.3108, 49.85345, 47.48175, 45.60637, 44.19613,
    43.44976, 43.47792,
  69.15096, 67.05114, 61.98462, 59.92418, 61.17197, 61.44666, 61.91141,
    62.0575, 62.33562, 62.28962, 61.4436, 60.12368, 58.87833, 57.79116,
    56.76159, 56.0521, 55.4526, 54.99775, 54.55376, 53.68206, 52.66772,
    52.26008, 52.69664, 51.7107, 51.13874, 48.53397, 46.36506, 44.73403,
    43.67178, 43.47039,
  67.76934, 65.93236, 61.15846, 59.04432, 60.45066, 61.01835, 61.90819,
    62.77128, 64.12942, 65.19621, 65.37022, 64.99767, 64.06007, 62.88829,
    61.54042, 60.50584, 59.61741, 58.63012, 57.46862, 56.21552, 54.74328,
    53.40047, 53.38383, 52.42598, 52.14383, 50.40339, 47.65692, 45.64222,
    44.37099, 43.64104,
  66.05016, 63.65543, 59.79351, 57.80801, 58.88908, 59.42578, 60.57312,
    62.29848, 64.57052, 66.27775, 67.42219, 68.68874, 69.88231, 69.66077,
    67.94863, 66.86921, 65.41461, 63.82281, 62.13564, 60.45078, 58.91332,
    57.00146, 54.83096, 53.98483, 53.64252, 52.66328, 50.32739, 46.75381,
    45.19218, 44.25232,
  64.46008, 61.53495, 56.94656, 55.17025, 55.83954, 56.39755, 58.16866,
    60.74701, 63.55778, 64.31488, 65.20353, 66.97767, 69.12051, 69.6565,
    68.42008, 67.44961, 66.31392, 64.8702, 63.15464, 61.89841, 60.15034,
    58.0836, 55.78586, 54.49316, 54.14882, 53.1457, 51.84308, 47.83545,
    45.44447, 44.62902,
  63.52562, 60.05237, 56.34918, 53.83702, 54.30439, 54.35989, 55.93904,
    58.7338, 61.08686, 61.60341, 62.87842, 64.90665, 67.13103, 67.90586,
    67.19269, 66.37917, 65.48688, 64.04429, 62.90159, 61.86753, 60.1101,
    58.38353, 56.12281, 54.84614, 54.50192, 53.26049, 51.97496, 49.22716,
    45.39553, 44.40901,
  62.05047, 59.23023, 55.72095, 53.3061, 53.62935, 53.24559, 54.05267,
    55.64265, 57.14389, 57.70893, 59.09853, 60.88021, 63.36531, 64.60329,
    63.85562, 63.70526, 63.09363, 62.1486, 61.01449, 60.4725, 59.09839,
    57.68215, 55.90369, 54.99997, 54.68552, 53.67825, 52.47781, 50.68967,
    46.91121, 44.25146,
  58.42665, 56.73624, 54.0077, 52.12334, 52.66934, 52.71272, 52.81432,
    53.54957, 53.97334, 53.85856, 54.17557, 55.297, 57.08699, 58.36938,
    58.46855, 58.38342, 58.09782, 57.59769, 57.32529, 57.12183, 56.68966,
    55.62237, 53.72454, 52.76792, 52.99895, 52.38267, 51.64982, 50.41451,
    48.38508, 45.23186,
  49.95488, 49.96395, 49.95839, 50.16784, 50.52466, 50.99793, 51.26022,
    50.99054, 50.04248, 50.12239, 49.81502, 49.48386, 49.83928, 50.47777,
    50.44255, 50.41109, 49.87498, 49.09908, 48.62059, 48.68507, 48.94457,
    49.73231, 49.61697, 48.95638, 49.02474, 48.83059, 48.18218, 46.81453,
    45.79185, 44.92239,
  47.69521, 48.05969, 48.37968, 48.18058, 48.8788, 50.24171, 50.6101,
    48.09197, 46.89886, 47.21313, 47.46396, 47.56813, 47.47075, 47.19823,
    46.76023, 46.63794, 45.85585, 44.8758, 44.75893, 44.67359, 44.63795,
    45.25558, 46.17783, 46.50434, 46.3277, 46.40744, 46.14471, 45.19804,
    44.26616, 43.58877,
  50.81348, 50.67147, 50.74086, 50.7773, 50.74026, 50.74502, 50.72093,
    50.71984, 50.79279, 50.90895, 51.11551, 51.30032, 51.32924, 51.58334,
    51.75219, 51.84946, 51.98843, 52.16122, 52.29902, 52.48961, 52.59034,
    52.44209, 52.38736, 52.53351, 52.67152, 52.18113, 51.81873, 51.88188,
    50.59545, 49.04145,
  50.94258, 50.88213, 50.94166, 50.9708, 50.93317, 50.88562, 50.86534,
    50.85603, 50.91455, 50.92632, 51.09911, 51.39382, 51.66232, 51.82004,
    51.91559, 52.15242, 52.35609, 52.69763, 53.11227, 53.50623, 53.81556,
    53.85349, 53.72878, 53.87527, 53.88699, 52.55001, 51.17703, 51.40455,
    50.36917, 49.22145,
  51.11377, 51.09341, 51.20785, 51.25497, 51.20239, 51.19485, 51.24044,
    51.30173, 51.37804, 51.40247, 51.45139, 51.65973, 51.86692, 51.98925,
    52.07588, 52.00418, 52.1476, 52.57552, 53.16249, 53.8485, 54.70156,
    55.38963, 55.50471, 55.37254, 54.79549, 53.2835, 52.00075, 51.28936,
    49.76651, 49.36004,
  51.25936, 51.24946, 51.43194, 51.4835, 51.42759, 51.47289, 51.57511,
    51.67281, 51.79467, 51.8121, 51.97375, 52.40233, 52.5875, 52.46841,
    52.53748, 52.50542, 52.34188, 52.41527, 53.00094, 53.78141, 54.5585,
    54.808, 54.9127, 55.33822, 54.79214, 53.88901, 53.15118, 52.44605,
    51.9209, 50.51097,
  51.31862, 51.34885, 51.57296, 51.63875, 51.56592, 51.67358, 51.893,
    51.91403, 51.8756, 51.84053, 52.1439, 52.91031, 53.5347, 53.56814,
    53.56749, 53.69342, 53.42104, 52.99108, 53.26432, 53.89864, 54.00479,
    53.53791, 53.84074, 54.39757, 54.51525, 54.10971, 53.91107, 54.50138,
    54.13172, 52.47134,
  51.16499, 51.31898, 51.66271, 51.80445, 51.70314, 52.06114, 52.75616,
    52.8611, 52.57598, 52.33802, 52.45451, 53.2808, 54.19226, 54.17803,
    54.51616, 54.98054, 54.56752, 53.8056, 53.46746, 53.77285, 53.61013,
    53.25886, 53.80181, 54.00274, 54.08191, 54.20716, 54.41463, 55.05383,
    54.04387, 51.67969,
  51.06709, 51.18183, 51.4629, 51.54885, 51.65633, 52.22673, 53.18574,
    53.71253, 53.68167, 53.3591, 53.15351, 52.73021, 52.14195, 52.4278,
    52.67846, 52.98222, 52.98212, 52.36547, 52.22636, 52.74692, 53.08288,
    53.43687, 53.88422, 54.21197, 54.14341, 54.01143, 54.50248, 54.56874,
    52.7922, 48.02847,
  51.43467, 51.26899, 51.44572, 51.46814, 51.48457, 52.12209, 52.77781,
    52.11933, 51.80278, 52.02499, 52.09512, 52.23672, 52.48923, 52.72918,
    52.92166, 53.12302, 53.06245, 52.80031, 52.48692, 52.55476, 52.99762,
    53.51239, 53.99259, 54.20862, 54.07328, 54.32024, 54.75825, 54.06812,
    52.15445, 48.22312,
  52.99155, 52.48199, 52.20548, 51.97156, 51.79668, 51.73905, 51.11681,
    51.38153, 51.7063, 51.88271, 52.10164, 52.32785, 52.6204, 53.3224,
    53.80073, 53.56837, 53.81707, 54.14878, 54.10969, 53.65119, 53.59291,
    53.88837, 53.99609, 53.72192, 53.78395, 54.46024, 54.28249, 52.96996,
    48.5334, 48.82845,
  55.8881, 55.44485, 54.60957, 53.94495, 53.46467, 52.30709, 50.85582,
    51.39299, 51.59481, 51.84439, 51.91616, 51.9455, 51.89993, 52.07852,
    52.27965, 52.97434, 53.64074, 54.10719, 54.28527, 54.42093, 54.76173,
    54.32981, 53.52678, 52.89153, 53.42415, 53.99396, 53.20832, 51.61517,
    48.29033, 48.23177,
  59.69166, 58.81292, 59.63995, 57.75192, 57.07961, 54.64391, 53.1059,
    52.25121, 52.18916, 52.74707, 51.97797, 50.89513, 50.83579, 51.04269,
    51.14977, 51.56139, 52.12945, 52.6369, 53.11387, 53.6479, 54.55929,
    54.39458, 53.35014, 53.16737, 53.52864, 53.02076, 51.62096, 48.56402,
    49.24523, 48.33358,
  64.0719, 62.54289, 64.37835, 64.66936, 62.27189, 59.007, 56.15537,
    53.27242, 51.75116, 52.41062, 52.02984, 51.54356, 51.71873, 51.78033,
    51.49191, 51.4655, 51.84895, 52.29387, 52.65393, 53.05674, 53.98016,
    54.00587, 53.2067, 53.54144, 53.72058, 52.46539, 49.01413, 51.5325,
    49.93301, 48.92449,
  56.90316, 58.46441, 60.1428, 61.88715, 62.91227, 61.43159, 55.4079,
    52.15166, 53.91275, 52.98194, 52.90826, 52.51802, 52.78065, 52.94004,
    52.56945, 51.53362, 52.01398, 52.49797, 52.83093, 53.13741, 53.74339,
    53.79892, 53.04584, 52.30756, 52.09043, 51.61077, 49.67085, 51.38225,
    50.87217, 49.56121,
  52.0876, 52.01149, 52.17074, 51.52268, 51.57293, 52.33255, 53.58214,
    53.99358, 52.59163, 53.01434, 53.39482, 52.9491, 52.97284, 53.19577,
    52.69836, 51.98019, 51.93628, 52.80574, 53.52506, 53.3397, 53.32537,
    53.00394, 52.04107, 51.52689, 49.23118, 49.59457, 49.17324, 48.70783,
    49.0158, 48.96048,
  53.93547, 53.92139, 53.46561, 52.7642, 52.32361, 52.43047, 53.10242,
    53.21875, 52.54912, 52.39616, 52.29139, 52.16262, 52.46153, 52.5633,
    52.38678, 52.39023, 51.97113, 52.43717, 53.048, 53.0316, 52.27726,
    51.94113, 51.12873, 49.99746, 50.88401, 50.28495, 49.46676, 48.8062,
    48.47586, 48.41753,
  52.79258, 53.21989, 53.39145, 53.21709, 53.13342, 53.55603, 54.02598,
    54.06837, 53.47434, 52.81704, 52.69815, 52.46618, 52.472, 52.89373,
    52.3082, 51.76173, 52.02302, 52.18959, 52.33936, 52.09356, 51.72463,
    51.41821, 50.6773, 49.86043, 50.34055, 50.18436, 49.33816, 48.84883,
    48.54693, 48.44691,
  52.77263, 52.49886, 52.53133, 52.5679, 52.60604, 52.59433, 53.18555,
    53.95717, 54.04544, 53.81286, 53.59787, 54.16068, 54.9631, 54.64981,
    53.7527, 53.27901, 53.20169, 53.29629, 53.03218, 52.31489, 51.69777,
    51.70789, 51.19539, 50.31036, 50.36012, 50.29256, 49.30736, 48.52417,
    48.42202, 48.40554,
  56.40845, 54.5128, 53.15214, 52.58748, 52.50443, 52.45069, 52.74517,
    53.25198, 53.65888, 53.70325, 54.27849, 55.0523, 55.43585, 55.54257,
    55.43099, 55.62836, 56.1245, 56.5225, 56.09566, 54.6418, 53.04847,
    52.45277, 52.07367, 51.46461, 50.66376, 50.11239, 49.32977, 48.38124,
    48.31916, 48.31238,
  66.1298, 61.54097, 56.22006, 52.87663, 53.28835, 52.74199, 52.89576,
    53.05567, 52.92825, 53.12872, 53.58171, 53.66377, 53.4875, 53.70004,
    53.86863, 54.82732, 56.51754, 58.28999, 58.89001, 57.95108, 56.09155,
    54.18948, 53.3055, 53.11214, 51.6659, 50.65244, 49.67626, 48.52372,
    48.29068, 48.33419,
  66.9537, 63.00388, 57.86633, 54.64791, 54.86097, 54.33187, 54.11486,
    53.85408, 53.72488, 53.83591, 53.76414, 53.3118, 53.19908, 52.74106,
    52.42586, 52.56912, 53.57129, 55.12268, 56.17076, 56.34702, 55.81266,
    54.83437, 53.93301, 53.54758, 52.9923, 51.3083, 50.09661, 48.71111,
    48.32886, 48.38956,
  68.45293, 65.28621, 59.95961, 57.1541, 57.38178, 56.86879, 56.5288,
    56.10418, 55.76341, 55.39946, 54.84353, 54.31182, 54.23265, 53.93659,
    53.55008, 53.49791, 53.82236, 54.47026, 54.96289, 54.7869, 54.60274,
    54.43807, 54.07679, 53.68213, 53.17078, 51.88368, 50.10297, 48.79266,
    48.28584, 48.35853,
  68.64585, 66.79869, 61.7949, 59.45962, 60.10336, 59.81805, 59.73998,
    59.48633, 59.33207, 58.95927, 58.03844, 57.11971, 56.49535, 55.89592,
    55.43137, 55.19514, 55.08395, 55.20523, 55.30965, 55.366, 55.30582,
    54.69218, 54.23064, 53.95115, 53.47251, 52.59199, 50.54758, 49.30964,
    48.45335, 48.31908,
  68.2326, 66.71312, 62.15763, 60.25113, 61.3456, 61.58464, 61.98301,
    62.37357, 63.23886, 63.53673, 63.06899, 62.70863, 61.96658, 61.04237,
    59.98282, 59.19556, 58.45401, 57.92982, 57.48043, 56.88442, 56.41702,
    55.57324, 54.68967, 54.37129, 54.12801, 53.15629, 51.84025, 50.31902,
    49.22449, 48.47746,
  66.95654, 65.10364, 61.30004, 59.74814, 60.4254, 60.64759, 61.62089,
    63.24976, 65.51727, 66.71365, 67.1243, 68.08355, 69.07971, 68.68305,
    67.09219, 65.75771, 64.32767, 63.04486, 61.89709, 60.62856, 59.23833,
    57.80773, 56.37791, 55.75347, 55.43675, 54.65327, 53.27232, 51.51611,
    50.34254, 49.11234,
  65.58485, 62.69191, 58.7704, 57.12763, 57.54852, 57.95227, 59.68589,
    62.50517, 65.3779, 65.72922, 65.9097, 67.24308, 68.96246, 69.3485,
    68.18379, 67.06243, 65.47884, 64.27431, 63.39402, 62.28255, 60.62045,
    58.81526, 57.142, 56.17591, 56.07715, 55.28882, 54.07339, 52.2645,
    50.78859, 49.69269,
  64.15102, 61.23496, 57.74437, 55.69569, 55.78261, 55.85437, 57.72486,
    60.87567, 63.32212, 63.46443, 64.31156, 65.74684, 67.6139, 68.40177,
    67.60368, 66.90436, 65.53513, 64.14864, 63.5721, 62.67761, 61.09689,
    59.51725, 57.88146, 56.87445, 56.54364, 55.52418, 54.40246, 52.65682,
    50.45702, 49.29667,
  62.11533, 59.73489, 56.72022, 54.42287, 54.6693, 54.31908, 55.46029,
    57.55302, 59.33889, 59.81601, 60.81491, 62.46006, 64.7383, 65.69168,
    65.34874, 65.07681, 64.29843, 63.26757, 62.71659, 62.08348, 60.76691,
    59.47254, 58.17897, 57.39989, 57.04071, 56.0923, 55.05146, 53.49224,
    51.78262, 49.08359,
  58.93078, 57.25691, 54.85587, 53.47699, 53.99125, 54.0176, 54.27331,
    55.1302, 55.70036, 55.83054, 56.21836, 57.37578, 59.33876, 60.46027,
    60.30481, 60.41083, 60.19378, 59.83533, 59.79508, 59.77839, 59.21946,
    58.05273, 56.73605, 56.1939, 55.97284, 55.24662, 54.45752, 53.51937,
    52.66066, 50.508,
  51.46493, 51.45044, 51.55285, 51.85447, 52.52677, 53.22934, 53.26915,
    53.0983, 53.26092, 53.23745, 53.00217, 52.73626, 52.71542, 52.95606,
    53.0883, 53.26973, 53.5278, 53.76389, 53.91411, 54.18672, 54.54329,
    54.97034, 54.88931, 54.28387, 53.98174, 53.66288, 53.20918, 52.12539,
    51.54109, 50.32335,
  51.62987, 51.41078, 51.44567, 51.43595, 52.00338, 52.82558, 53.18331,
    52.89398, 52.11992, 52.93079, 53.10382, 52.86457, 52.38163, 51.93921,
    51.71671, 51.79796, 51.44642, 50.29039, 50.29762, 50.24866, 50.14887,
    50.79412, 51.56132, 51.70391, 51.55311, 51.77775, 51.4167, 50.30107,
    49.34853, 48.50606,
  53.63323, 53.57953, 53.78809, 53.95079, 54.07856, 54.26609, 54.45444,
    54.66626, 54.93121, 55.31131, 55.81987, 56.09342, 55.98829, 56.44432,
    57.07995, 57.73581, 58.53491, 59.56781, 60.66754, 61.69193, 62.25546,
    62.24994, 62.37032, 62.78106, 63.08422, 62.62869, 62.77975, 62.87583,
    60.25805, 56.74828,
  52.95473, 52.95709, 53.08978, 53.27785, 53.27003, 53.34857, 53.5383,
    53.8127, 54.18164, 54.6224, 55.20396, 55.89191, 56.53119, 56.84108,
    57.35884, 58.24506, 58.99982, 60.11926, 61.37872, 62.50621, 63.1722,
    63.39291, 63.42456, 63.93755, 64.10506, 62.78102, 61.82969, 62.25787,
    60.19994, 57.5431,
  53.20069, 53.27349, 53.59034, 53.7529, 53.83839, 53.93213, 54.07046,
    54.34805, 54.6378, 54.95616, 55.42003, 56.04086, 56.74699, 57.61304,
    58.35199, 58.7163, 59.50418, 60.64147, 61.80426, 63.18169, 64.56911,
    65.42345, 65.61858, 65.74271, 65.22474, 63.44386, 62.28469, 61.77193,
    59.30418, 57.99673,
  53.39319, 53.48771, 53.87675, 54.15282, 54.37333, 54.67226, 54.98012,
    55.25882, 55.62389, 55.9432, 56.3009, 56.91644, 57.40612, 57.77284,
    58.70778, 59.48301, 59.68682, 59.96261, 61.31774, 62.94063, 64.58315,
    65.38702, 65.8034, 66.58356, 66.14143, 64.66988, 63.01028, 61.96489,
    61.43095, 58.18536,
  53.71039, 53.69023, 54.0381, 54.17079, 54.27924, 54.53497, 55.0113,
    55.44146, 55.98111, 56.51069, 56.91832, 57.73833, 58.49207, 58.92785,
    59.52785, 60.33284, 60.52074, 60.17315, 61.03389, 62.60793, 63.63846,
    63.8509, 64.59206, 65.72665, 66.12888, 65.12344, 63.67315, 63.8703,
    63.58883, 61.9405,
  53.77169, 54.08873, 54.55454, 54.86296, 54.72508, 54.93278, 55.67393,
    55.92249, 55.8954, 56.16716, 56.89455, 58.07182, 59.28233, 59.69346,
    60.66949, 61.81713, 62.12631, 61.74072, 61.53765, 62.60547, 63.21159,
    63.41224, 64.3428, 65.0077, 65.32052, 65.02541, 64.34566, 64.98047,
    63.88692, 61.34417,
  53.62697, 54.03644, 54.63745, 55.03711, 55.13063, 55.6517, 56.64956,
    57.1246, 57.15566, 57.17034, 57.44649, 57.48714, 57.38884, 58.31156,
    59.40133, 60.59295, 61.29395, 61.0916, 61.016, 62.2658, 63.15724,
    63.91186, 64.61446, 65.34671, 65.24682, 64.43973, 64.63508, 64.46364,
    62.67717, 55.43053,
  53.95711, 54.26966, 54.94247, 55.3955, 55.57382, 56.44318, 57.32677,
    56.8123, 56.62201, 57.16409, 57.51676, 58.00794, 58.64997, 59.65067,
    60.56933, 61.45467, 62.23847, 62.41435, 62.19936, 62.77933, 63.63891,
    64.60262, 65.49054, 65.82083, 65.15617, 65.01151, 65.47188, 64.50365,
    62.30617, 56.2742,
  56.03628, 56.0838, 56.16597, 56.16928, 55.87055, 56.18368, 56.18283,
    57.00233, 57.99427, 58.75324, 59.35224, 59.87139, 60.66769, 62.50739,
    63.75821, 63.05475, 63.82806, 64.87704, 65.0645, 64.57227, 64.7054,
    65.74747, 66.58994, 66.0456, 65.15141, 65.88045, 65.06493, 63.1828,
    57.62203, 56.6684,
  58.42081, 59.12194, 58.57983, 58.62233, 58.02472, 56.68014, 55.47502,
    56.50597, 57.09505, 58.34332, 59.59874, 60.63984, 60.90031, 61.08192,
    61.34836, 62.986, 64.0654, 64.69056, 65.15424, 65.92554, 66.92589,
    66.28511, 65.09292, 63.51382, 64.00543, 64.70044, 63.50907, 61.46995,
    55.99029, 54.97955,
  58.84546, 58.47595, 59.94424, 59.13916, 60.0357, 58.76631, 57.91215,
    57.55866, 58.10513, 59.13424, 58.58728, 57.30047, 57.82081, 58.47985,
    59.18618, 59.98546, 61.00295, 61.80119, 62.62822, 63.91938, 66.077,
    65.8127, 63.51227, 62.66435, 62.9529, 62.5318, 61.14368, 56.26328,
    56.64835, 55.19957,
  63.53364, 61.30288, 63.36252, 64.50452, 63.22897, 61.69836, 60.22688,
    57.9074, 56.33054, 57.07156, 57.27274, 57.32373, 58.33343, 59.32914,
    59.42883, 59.74653, 60.30961, 61.06052, 61.8419, 62.9428, 64.80731,
    65.01839, 63.20124, 63.59917, 63.38422, 61.94654, 56.80343, 60.74857,
    57.66664, 56.14572,
  62.4445, 63.61597, 65.14919, 66.66153, 67.09314, 65.63902, 60.09093,
    57.40491, 59.34529, 58.38609, 58.68192, 58.57653, 59.90594, 60.88849,
    60.38734, 59.90397, 60.62491, 61.3569, 62.10283, 63.35348, 64.38564,
    64.16788, 63.11003, 62.285, 61.95085, 61.23294, 58.15613, 59.72854,
    59.1807, 57.24177,
  56.32826, 57.08726, 56.95935, 56.5777, 56.98243, 57.92548, 59.37411,
    59.81572, 58.50357, 59.19004, 60.11893, 60.00246, 61.25163, 61.85921,
    61.23992, 60.46779, 60.54107, 61.78044, 63.00883, 63.39213, 63.27068,
    62.84522, 61.99281, 61.36459, 58.68424, 58.26593, 57.01494, 56.36548,
    56.89431, 56.59471,
  56.46244, 56.92672, 56.91836, 56.72586, 56.97443, 58.54326, 60.53617,
    59.80478, 58.70865, 58.78764, 58.73484, 58.88805, 59.85468, 60.80644,
    60.96167, 60.43183, 60.44644, 61.49569, 63.19244, 63.62686, 62.09729,
    61.96327, 60.97853, 59.78594, 60.17351, 58.77589, 57.27394, 56.31937,
    55.7746, 55.54291,
  56.4844, 57.16857, 57.4895, 57.38058, 57.44886, 58.39393, 59.58034,
    59.67614, 59.0359, 58.7583, 59.14934, 58.88139, 58.96767, 60.02997,
    59.90081, 59.81187, 60.42079, 61.116, 62.30825, 62.38865, 61.48506,
    61.55782, 60.49747, 59.22848, 59.70009, 58.92529, 57.03409, 56.43584,
    55.9296, 55.62105,
  55.04525, 55.07585, 55.5971, 56.1158, 56.73284, 57.27945, 58.25293,
    59.40788, 59.78694, 59.65185, 59.30696, 60.52301, 62.04585, 61.39952,
    60.37873, 60.06316, 60.2448, 60.99024, 62.0339, 61.89355, 60.94228,
    61.58706, 60.9695, 59.6576, 59.34673, 59.19597, 57.03374, 55.59776,
    55.6244, 55.51142,
  56.10526, 55.40485, 54.96624, 55.24524, 55.76807, 56.44238, 57.3385,
    58.49564, 59.38529, 59.75623, 61.23188, 62.82745, 63.30087, 63.71075,
    63.34707, 62.85312, 62.92633, 63.80204, 64.51849, 63.4897, 61.68891,
    61.87772, 61.66878, 61.151, 58.94086, 57.86349, 57.01871, 55.29141,
    55.27918, 55.22008,
  64.15202, 60.57851, 56.30052, 53.87337, 54.87043, 55.08669, 55.96672,
    56.96973, 57.6759, 58.65862, 60.0852, 60.68567, 60.62497, 61.83501,
    62.60868, 63.86527, 66.22043, 68.76649, 69.54095, 68.23601, 65.50702,
    63.76295, 62.97263, 62.26416, 59.45203, 57.77348, 56.93337, 55.66615,
    55.25556, 55.22369,
  64.1421, 60.62561, 56.49885, 54.02813, 54.6932, 54.7748, 55.3164, 55.96132,
    56.83563, 58.05649, 58.57156, 57.96249, 58.7295, 59.27304, 59.74186,
    60.40111, 62.10701, 64.61604, 66.57909, 67.24516, 66.5324, 65.17197,
    63.89314, 63.17017, 61.56754, 58.65795, 57.28225, 55.89268, 55.22311,
    55.23312,
  65.1573, 61.96008, 57.61722, 55.34834, 55.61683, 55.49183, 55.67821,
    56.04199, 56.69886, 57.29968, 57.04416, 56.70863, 57.68142, 58.1145,
    58.34476, 58.89709, 60.21671, 61.94998, 63.66879, 64.53429, 65.12682,
    65.48982, 64.91461, 63.88826, 62.77861, 59.70835, 57.15716, 55.83651,
    55.20047, 55.23106,
  67.25945, 64.80457, 60.40916, 58.23707, 58.66202, 58.23707, 58.23984,
    58.24098, 58.77921, 58.97865, 58.13515, 57.8204, 58.28534, 58.49792,
    58.74113, 59.33319, 60.12882, 61.30243, 62.57916, 63.75527, 64.90419,
    65.24709, 65.21043, 64.88062, 63.84682, 61.39004, 57.79983, 56.6575,
    55.43256, 55.18053,
  69.12572, 67.61961, 63.35585, 61.51124, 62.52811, 62.64613, 62.60076,
    62.52727, 63.158, 63.13671, 62.32361, 62.58613, 62.67364, 62.61198,
    62.43151, 62.62658, 62.91821, 63.09291, 63.58496, 64.2866, 65.07823,
    65.10782, 64.61161, 64.71519, 64.85797, 63.30607, 60.35267, 58.57235,
    56.84351, 55.39374,
  69.59908, 68.09541, 64.83399, 63.3684, 63.97863, 64.13158, 65.08831,
    66.34897, 68.4693, 68.85844, 68.35232, 69.49753, 70.71947, 70.99216,
    70.32006, 69.85509, 69.26964, 68.63907, 67.84805, 67.63062, 67.67838,
    67.1129, 66.0528, 65.61886, 65.69896, 65.21672, 63.45176, 60.87721,
    59.01356, 56.49105,
  69.5285, 66.4419, 62.75418, 61.18965, 61.73468, 62.27697, 64.06986,
    66.93302, 69.88792, 69.56352, 69.02155, 70.55526, 72.08942, 72.70412,
    72.19636, 71.81154, 71.21647, 70.7564, 70.2261, 69.90597, 69.37975,
    68.40036, 67.04414, 66.1648, 66.24811, 65.83788, 64.66994, 62.51202,
    60.84562, 58.17937,
  69.01856, 66.4503, 63.03481, 60.94378, 61.02676, 61.36081, 63.67038,
    67.06361, 69.09133, 68.43704, 69.04691, 70.45996, 72.31134, 72.93059,
    72.21669, 72.08258, 71.71121, 71.43974, 71.38554, 71.27765, 70.91127,
    69.92359, 68.38756, 67.38096, 67.15153, 66.34348, 65.357, 63.22687,
    59.75714, 57.31154,
  67.07069, 64.60316, 61.8895, 60.01108, 60.22064, 60.15078, 61.89217,
    64.08299, 65.30782, 65.64167, 67.01246, 68.72601, 70.62231, 71.4406,
    71.14446, 71.11064, 71.01675, 71.01711, 71.13512, 71.47495, 71.18732,
    70.95206, 69.9633, 68.993, 68.61764, 67.86008, 67.0197, 65.11618, 61.848,
    56.21764,
  63.48388, 61.80528, 60.06541, 59.32763, 60.2463, 60.29685, 60.66004,
    61.17572, 61.23173, 61.84671, 62.86214, 64.53056, 66.59393, 67.74123,
    67.83115, 67.89509, 68.11802, 68.30892, 69.02877, 69.85471, 69.59932,
    68.69697, 67.35059, 66.79947, 66.8874, 66.43015, 65.77941, 65.42891,
    64.16643, 60.03193,
  56.41262, 56.40261, 56.81515, 57.56746, 59.19481, 60.82318, 60.48391,
    59.52272, 59.57566, 59.93923, 60.02179, 60.27324, 60.6921, 61.38342,
    61.89722, 62.38118, 62.89364, 63.43586, 63.70671, 63.99831, 64.59152,
    64.97397, 64.70403, 63.99965, 63.96655, 63.89852, 63.3545, 62.43426,
    62.24198, 60.31823,
  58.10649, 58.09336, 58.43943, 58.77168, 60.24081, 62.30419, 63.22976,
    61.99684, 61.59895, 62.25829, 62.80701, 63.09227, 62.85744, 62.33116,
    61.93605, 61.8428, 61.50973, 60.61381, 60.59576, 59.99491, 58.87168,
    59.64954, 60.13266, 60.33172, 60.68693, 61.60135, 61.63137, 59.39582,
    57.12087, 55.29485,
  55.77842, 56.12904, 56.39168, 56.80653, 56.92738, 57.19562, 57.62163,
    58.10773, 58.29819, 58.49585, 58.94262, 58.90065, 57.8343, 57.88104,
    57.76283, 57.13128, 57.04718, 57.21365, 57.36283, 57.74565, 57.83933,
    57.44685, 57.57521, 58.27737, 58.83996, 58.60229, 59.72523, 60.02762,
    56.71994, 52.398,
  58.14888, 58.45198, 58.52228, 58.94886, 58.92496, 58.93325, 59.18339,
    59.38914, 59.52474, 59.65631, 59.91307, 60.2506, 60.24653, 59.40279,
    58.72829, 58.51558, 57.91224, 57.90236, 58.14, 58.35595, 58.185,
    57.90105, 57.8991, 58.65809, 59.01863, 58.17627, 58.52705, 59.62021,
    57.15843, 53.86104,
  58.03559, 58.43162, 58.94593, 59.4176, 59.77457, 59.9635, 60.04379,
    60.16202, 60.2482, 60.25877, 60.25374, 60.322, 60.38757, 60.47215,
    60.2482, 59.25422, 58.77163, 58.807, 58.85728, 58.97625, 59.29308,
    59.56703, 59.79342, 60.26025, 60.14067, 58.96767, 58.80856, 58.89962,
    57.10737, 55.07626,
  59.29556, 59.65958, 60.23175, 60.71251, 61.14455, 61.58281, 61.60255,
    61.43676, 61.37806, 61.2005, 61.02399, 61.23463, 61.06014, 60.37105,
    60.74589, 60.91555, 59.71169, 58.59386, 58.9971, 59.47256, 59.99235,
    60.22187, 60.75806, 61.9088, 62.20602, 61.18276, 59.17891, 57.79743,
    57.11478, 53.52368,
  59.9875, 59.96252, 60.52511, 60.87515, 61.07984, 61.28376, 61.48653,
    61.40948, 61.22961, 60.9024, 60.79439, 61.44441, 61.72716, 61.58054,
    61.47594, 61.59737, 60.71761, 58.92951, 58.91987, 59.50919, 59.48207,
    59.15913, 59.81568, 61.37439, 62.70071, 61.51528, 58.62415, 58.41265,
    58.38769, 56.97386,
  60.06135, 60.66425, 61.57576, 62.1919, 62.06956, 62.49164, 63.33502,
    63.11436, 62.43691, 62.068, 62.08637, 62.65343, 63.20088, 62.67282,
    62.93753, 63.60905, 62.60646, 60.48495, 58.76242, 59.13878, 59.03916,
    58.76999, 59.36483, 60.54944, 61.70731, 60.98646, 58.86491, 59.36707,
    58.90872, 56.98912,
  60.47047, 61.11826, 61.90072, 62.36142, 62.16846, 62.36549, 62.74842,
    62.46394, 61.8741, 61.61809, 61.64248, 61.67598, 61.61057, 62.1925,
    62.50454, 62.6104, 62.49269, 60.75212, 58.79017, 59.26489, 59.27798,
    59.46445, 60.15614, 61.51161, 61.48635, 59.67704, 59.33926, 59.17781,
    58.39281, 52.99806,
  61.27087, 61.99004, 62.79388, 63.29351, 62.91365, 62.99981, 63.61371,
    62.66348, 61.60559, 61.59218, 61.53616, 61.66045, 61.92233, 62.55735,
    63.0346, 63.39676, 63.6916, 62.89835, 60.92444, 60.4914, 60.35392,
    60.86407, 62.00209, 62.56937, 61.34134, 60.36895, 60.7718, 60.17886,
    58.6825, 53.45703,
  63.63864, 64.17196, 64.79173, 64.7472, 63.64802, 63.68383, 63.96959,
    64.45485, 65.12116, 65.61522, 66.06116, 66.32529, 66.80157, 69.35135,
    70.89967, 67.89622, 67.93823, 68.25451, 67.10258, 64.59831, 63.0842,
    64.3126, 66.11214, 65.02615, 62.42131, 63.16774, 61.79655, 59.63076,
    57.17382, 52.62052,
  69.59818, 71.51913, 71.17124, 71.71736, 69.62173, 67.4284, 65.74121,
    66.39278, 66.78778, 68.83705, 70.2755, 71.07931, 70.29403, 68.50859,
    66.7391, 68.26926, 68.96329, 68.87033, 68.6587, 68.59267, 67.87029,
    66.25712, 64.41948, 61.67704, 61.03473, 60.97442, 59.88752, 57.49342,
    52.27276, 49.84462,
  67.21131, 67.04551, 68.83691, 68.80677, 69.43818, 68.0533, 66.81059,
    66.33199, 66.79604, 66.80325, 64.83578, 60.78614, 60.18663, 60.1134,
    60.37535, 60.93337, 61.73062, 62.24257, 62.87961, 63.51082, 64.69799,
    63.86702, 59.50354, 57.73424, 57.88826, 57.67358, 56.67046, 52.47398,
    51.85526, 50.02908,
  71.33031, 69.13454, 72.3913, 73.10833, 71.12258, 68.89597, 66.61567,
    63.70894, 61.24747, 60.70285, 60.01667, 59.07589, 59.62978, 60.4592,
    60.43899, 60.4166, 60.59435, 61.31416, 62.7103, 64.15841, 64.3982,
    62.36708, 58.48911, 58.76058, 58.38269, 57.0193, 52.76811, 54.71033,
    53.11019, 51.14577,
  74.87846, 76.539, 78.48637, 78.60815, 77.09457, 73.67759, 66.43021,
    62.59562, 63.21679, 61.02846, 61.07405, 60.40092, 61.1758, 61.88817,
    61.37478, 60.49257, 60.80759, 61.25793, 62.79737, 65.39142, 64.03708,
    60.56067, 58.94542, 57.92152, 57.80207, 57.00173, 53.87541, 54.70012,
    54.81923, 52.33995,
  67.87579, 68.6737, 69.10742, 67.94573, 67.29005, 68.33143, 70.04485,
    69.65875, 65.76659, 64.91851, 64.53379, 62.29728, 63.37202, 63.99994,
    62.17464, 60.80169, 60.5304, 60.75357, 61.3694, 61.7541, 60.72906,
    59.17645, 58.09781, 57.20359, 56.43356, 55.10287, 52.66585, 52.00157,
    52.51962, 51.78791,
  65.01899, 66.02287, 66.58228, 66.59364, 66.12523, 66.83749, 69.94267,
    69.93392, 66.09934, 64.68417, 63.36587, 62.59595, 63.29376, 63.53662,
    62.6874, 61.87544, 61.23946, 61.97089, 63.29317, 62.80447, 58.64171,
    58.40286, 57.20627, 56.74887, 56.9804, 54.87491, 52.98329, 51.81538,
    51.24508, 50.6161,
  66.27102, 67.2215, 67.9134, 67.35149, 66.28717, 67.18365, 68.54722,
    67.53575, 65.29555, 63.69972, 63.62882, 62.18243, 61.43799, 62.83634,
    62.00212, 61.3395, 61.59372, 61.59167, 62.23999, 61.12457, 58.17748,
    57.89631, 56.61186, 56.55321, 57.00016, 54.79739, 53.01745, 51.89417,
    51.38066, 50.68693,
  64.70272, 64.46308, 64.93685, 65.44324, 65.59302, 65.10364, 65.87035,
    66.98425, 66.31137, 65.15701, 63.19619, 64.15422, 66.63912, 64.67333,
    62.2458, 61.61366, 61.16784, 61.34084, 62.25516, 61.21016, 57.63711,
    58.00545, 57.00975, 56.68471, 56.91681, 55.40306, 52.75483, 50.74522,
    50.73074, 50.46405,
  64.17673, 64.64957, 64.72074, 65.41468, 66.03696, 66.44025, 66.12885,
    65.79853, 65.36856, 64.72261, 66.30173, 69.00033, 68.58321, 65.85142,
    64.87191, 63.46929, 62.06432, 62.60273, 63.82574, 61.20463, 57.85762,
    57.50055, 57.03732, 56.8891, 54.89671, 53.44994, 52.64381, 50.32001,
    50.26512, 50.05935,
  68.90864, 67.18504, 64.69894, 63.09303, 63.5588, 63.20315, 63.32959,
    63.65541, 63.21893, 63.6, 64.67975, 64.26541, 62.37266, 62.81313,
    62.54617, 63.48465, 65.58835, 67.88913, 68.74519, 66.16868, 61.25975,
    58.72454, 57.78719, 57.45974, 54.48128, 52.57972, 51.98399, 50.63836,
    50.22303, 50.08237,
  68.53143, 66.89847, 64.59394, 63.04609, 63.72403, 63.72796, 63.42891,
    63.27181, 63.78268, 65.57887, 66.15402, 63.88458, 63.30456, 62.57725,
    62.02713, 62.39946, 64.49998, 66.54425, 65.59225, 64.58604, 62.7209,
    60.3579, 58.60849, 58.07184, 56.6515, 53.35009, 51.99281, 50.65796,
    50.17401, 50.05767,
  68.57306, 67.512, 64.43372, 62.84646, 63.26269, 63.18597, 62.89209,
    62.82773, 63.57335, 64.70045, 64.02522, 62.6033, 63.10284, 62.5248,
    61.66496, 60.90443, 61.00809, 61.06401, 61.28387, 61.13678, 60.81747,
    61.13024, 60.04005, 59.03708, 57.89318, 54.16076, 51.60057, 50.72364,
    50.16686, 50.0905,
  68.6583, 66.9707, 64.57339, 63.08128, 63.17469, 62.64077, 62.70216,
    62.85738, 63.81622, 63.99765, 61.89624, 60.56149, 61.06391, 61.10837,
    60.87599, 60.85302, 60.70236, 60.69341, 60.91549, 60.73728, 60.37272,
    60.26807, 60.52655, 60.37581, 58.888, 55.82231, 52.03952, 51.31482,
    50.433, 50.0797,
  70.31672, 69.74779, 66.22044, 64.84313, 65.41086, 65.02288, 64.72559,
    64.27341, 65.0666, 64.75243, 62.51298, 62.08931, 62.43477, 62.26203,
    61.36287, 61.65776, 61.44873, 60.62964, 60.22421, 59.81961, 59.29153,
    59.05477, 58.78444, 59.24647, 59.75953, 58.22479, 54.65661, 53.47824,
    52.11086, 50.29533,
  70.73873, 70.23122, 68.36274, 66.56889, 66.66959, 66.06377, 66.55435,
    67.58944, 69.49848, 68.81828, 66.50636, 66.31734, 67.09914, 67.36857,
    65.96213, 65.8363, 65.39909, 64.47889, 63.07318, 62.09939, 60.89405,
    59.93256, 59.31153, 59.11968, 59.68974, 60.18686, 58.67443, 55.34306,
    54.07338, 51.28371,
  73.09481, 71.31358, 67.56458, 65.71829, 65.71865, 65.51845, 66.12271,
    68.12547, 70.94419, 70.25883, 67.39974, 67.21674, 67.61617, 68.00161,
    67.92692, 68.1018, 67.77612, 67.15587, 65.55256, 63.98914, 62.62244,
    61.69561, 60.76789, 60.14412, 60.19074, 60.61473, 60.37492, 58.19437,
    57.15005, 53.94481,
  74.00053, 72.61454, 69.55179, 66.8483, 65.96448, 65.57872, 67.41229,
    70.26566, 71.187, 69.71969, 68.55582, 68.07335, 68.73126, 68.89502,
    68.12143, 68.42824, 68.53551, 68.09332, 66.81927, 65.45854, 64.23543,
    63.26919, 61.92087, 61.10244, 61.22872, 60.83936, 60.53896, 58.89735,
    56.06153, 52.92629,
  73.6074, 72.03659, 69.46403, 67.12425, 66.80119, 65.9047, 67.5071,
    69.37789, 69.4764, 69.02053, 68.74437, 68.1423, 68.40507, 68.67577,
    68.59679, 68.66589, 68.85403, 68.8202, 67.7917, 66.44475, 65.51456,
    65.35772, 64.55287, 63.25271, 62.95679, 62.92544, 62.71614, 61.17669,
    57.38573, 50.87565,
  72.5423, 70.54289, 69.52696, 68.7095, 69.54066, 69.15911, 68.826, 68.43421,
    67.58037, 67.94917, 67.84419, 67.37178, 67.61932, 68.15836, 68.20184,
    68.10593, 67.89598, 67.61617, 67.27002, 66.9164, 65.56263, 64.23936,
    62.92714, 62.5294, 62.57123, 62.44113, 62.21763, 62.37978, 60.98128,
    56.45385,
  66.05772, 66.0284, 66.39272, 66.66515, 68.25438, 69.74189, 68.90002,
    66.17957, 65.19491, 65.23502, 65.06726, 65.23464, 64.88717, 64.46803,
    64.28572, 63.84835, 63.24194, 62.75591, 61.78811, 60.3346, 59.76129,
    59.46539, 58.77855, 58.15608, 58.69, 59.02511, 58.92327, 58.40903,
    58.512, 57.58202,
  65.09943, 65.56313, 65.48367, 64.05587, 65.28148, 67.45964, 67.77747,
    64.8914, 63.1026, 63.46474, 63.84072, 64.20879, 64.00117, 63.0197,
    61.70877, 61.01511, 59.59188, 58.4543, 58.1571, 57.75321, 55.67298,
    55.41302, 55.41573, 55.37947, 56.13591, 57.7301, 57.51455, 56.04501,
    52.80306, 50.14122,
  43.87959, 44.28608, 44.68357, 45.17487, 45.54947, 45.97269, 46.46381,
    47.04251, 47.70462, 48.52691, 50.24222, 50.52008, 48.67478, 49.26432,
    49.56209, 48.91503, 48.62687, 48.72065, 49.09573, 50.43613, 51.21382,
    50.53196, 51.21124, 52.54344, 53.2063, 52.69269, 55.56367, 55.88457,
    45.9853, 42.53747,
  51.52081, 52.36627, 52.4722, 53.70583, 54.02742, 54.45631, 55.37271,
    56.25546, 57.2942, 58.36782, 59.56429, 61.09058, 61.91363, 60.96573,
    60.13836, 59.98503, 57.9922, 57.36401, 57.63132, 58.09819, 57.78392,
    57.08875, 57.27872, 59.84103, 63.93672, 62.46407, 58.04416, 58.92632,
    47.32161, 43.799,
  57.04174, 58.04036, 58.88823, 59.28109, 59.33646, 59.43396, 59.57312,
    59.71214, 59.88409, 60.0089, 60.19527, 60.57493, 60.87604, 61.4016,
    62.1358, 62.88527, 64.31375, 65.94621, 67.07751, 67.63915, 67.85528,
    67.87267, 67.85013, 68.03863, 68.14124, 67.5088, 64.49269, 57.80844,
    47.59311, 44.97309,
  59.44825, 59.37859, 59.55045, 59.70373, 59.89025, 60.26638, 60.51474,
    60.63084, 60.87, 60.92552, 60.95597, 61.45543, 61.76414, 61.78148,
    62.83662, 64.26572, 65.18962, 66.23119, 67.69737, 68.43984, 68.83984,
    68.85744, 68.72286, 69.61222, 69.96818, 68.50401, 67.09495, 56.13518,
    47.77802, 43.46177,
  60.32186, 60.16117, 60.36712, 60.53016, 60.54471, 60.81959, 61.31998,
    61.55308, 61.76336, 61.75007, 61.74401, 62.22554, 62.62333, 62.93834,
    63.46812, 64.63717, 65.69525, 66.44728, 67.63091, 68.64261, 69.11467,
    68.65234, 68.65273, 69.05308, 69.58251, 68.57588, 65.74522, 65.07894,
    60.603, 47.46312,
  61.17544, 61.33518, 61.69478, 61.77163, 61.35535, 61.40757, 62.06813,
    62.20594, 61.94795, 61.89646, 62.12183, 62.8466, 63.56756, 63.54809,
    63.93023, 65.40907, 67.43228, 67.98759, 67.76495, 68.38382, 68.25561,
    66.83115, 67.69108, 68.14143, 68.5359, 67.66423, 66.1003, 66.83128,
    66.69955, 45.71258,
  62.18065, 62.29256, 62.47491, 62.3713, 61.80498, 61.75413, 62.25789,
    62.2926, 61.889, 61.78378, 61.90379, 61.99326, 62.0309, 62.30178,
    62.6384, 64.06406, 66.35927, 67.32426, 67.43077, 67.9495, 66.3338,
    64.68382, 65.35013, 67.70777, 67.32413, 63.36409, 66.50852, 66.89477,
    62.98811, 42.63865,
  62.56769, 62.52735, 62.54387, 62.36559, 61.67731, 61.48463, 61.7886,
    61.43003, 60.89478, 60.88864, 61.07467, 61.25629, 61.3743, 61.64933,
    62.32546, 64.01347, 66.33286, 67.81773, 67.72038, 66.21938, 64.97558,
    65.04382, 67.08733, 68.15691, 65.11436, 63.9157, 67.61897, 67.36373,
    53.1512, 43.07752,
  63.94732, 63.91786, 63.9462, 63.52466, 62.74908, 62.74356, 62.83592,
    63.27081, 63.92397, 64.19162, 64.46132, 64.76705, 65.08964, 66.57097,
    67.67085, 67.20222, 69.02721, 71.23405, 72.03387, 71.24238, 70.4251,
    70.89252, 71.72321, 70.8072, 68.83566, 68.85976, 68.16741, 60.97552,
    46.30984, 42.5406,
  70.73836, 71.15642, 70.75204, 70.86696, 69.63558, 67.71224, 66.93838,
    67.677, 68.1211, 68.98147, 69.70872, 70.57828, 70.38845, 69.43193,
    69.05084, 70.81346, 72.38382, 73.13439, 72.70366, 72.30274, 72.21561,
    71.18958, 69.91595, 68.10651, 68.09196, 69.25054, 67.31776, 47.56924,
    42.5809, 40.99634,
  71.83364, 72.00852, 73.76849, 73.73514, 74.90324, 73.73508, 72.32858,
    71.46513, 71.07755, 71.54063, 71.28857, 66.48615, 65.79822, 65.57256,
    66.27442, 67.78897, 69.62801, 70.50218, 70.37666, 70.02127, 70.51311,
    67.52489, 58.94209, 54.38897, 55.3257, 54.07969, 47.11133, 42.34992,
    41.84148, 40.94506,
  72.64429, 69.10458, 71.93108, 73.30376, 72.84196, 71.73319, 70.90694,
    68.18267, 65.24336, 64.76781, 63.92116, 62.82391, 62.99213, 63.3514,
    63.51426, 64.62187, 66.32977, 67.76056, 65.43184, 64.2589, 65.1858,
    60.76369, 52.91892, 58.10053, 60.63332, 47.72265, 42.16659, 42.87069,
    42.28019, 41.38791,
  77.1451, 76.97594, 78.2925, 78.98431, 77.96063, 75.07497, 68.72812,
    65.62797, 66.14038, 63.61074, 64.08851, 63.55871, 63.74324, 64.02401,
    63.59972, 64.07848, 66.17334, 67.77375, 67.42731, 68.31835, 66.26735,
    58.14175, 53.49495, 54.00673, 54.31071, 45.937, 42.99693, 43.20431,
    43.174, 41.98262,
  72.62904, 72.53851, 72.40456, 70.60238, 69.2458, 68.51126, 68.52164,
    69.13906, 66.95207, 66.69801, 67.40937, 65.83936, 67.14191, 67.64114,
    65.85651, 65.27766, 66.59977, 68.62152, 69.68837, 69.43339, 65.23032,
    58.07278, 57.31591, 49.13399, 45.07879, 44.14276, 42.76841, 42.20078,
    42.39902, 41.85263,
  65.80186, 65.35426, 65.10674, 64.72195, 64.81232, 66.01649, 69.54263,
    70.89809, 68.53049, 68.61527, 68.14436, 67.56999, 67.49509, 66.55316,
    65.53162, 65.03912, 66.28457, 68.21613, 69.90476, 69.42351, 59.44522,
    55.66795, 48.4871, 45.82684, 44.51638, 43.83571, 42.73296, 41.95018,
    41.62405, 41.27959,
  67.02335, 67.3055, 67.74538, 67.71587, 67.76739, 68.89554, 70.03865,
    69.78819, 69.36024, 68.71154, 68.0217, 66.01065, 64.93041, 65.28178,
    64.3232, 64.60854, 66.32372, 67.88776, 67.1046, 62.22106, 51.17485,
    49.92667, 46.83002, 45.57988, 44.72103, 43.71203, 42.64649, 42.03336,
    41.60228, 41.21239,
  67.20782, 66.98667, 67.06345, 67.22422, 67.75838, 67.80894, 68.33295,
    68.91413, 68.39879, 67.73193, 66.35266, 66.39532, 67.19962, 65.31358,
    64.18105, 64.54918, 66.2781, 67.43262, 66.71822, 63.58056, 49.9479,
    49.83984, 47.36704, 45.62844, 44.29638, 43.8035, 42.6009, 41.57735,
    41.37333, 41.1541,
  65.43026, 65.70445, 65.67501, 65.96877, 66.12072, 66.55243, 66.81425,
    67.20341, 67.53763, 66.72345, 66.91788, 67.29559, 66.24061, 65.30053,
    65.19724, 64.93885, 65.94186, 63.11683, 64.72047, 60.62488, 50.11508,
    48.90095, 46.73028, 45.26679, 43.33365, 42.82538, 42.32169, 41.26816,
    41.08319, 40.97255,
  67.51959, 66.14335, 64.75031, 64.07188, 64.59915, 64.70998, 65.12344,
    65.57658, 65.45157, 65.42017, 65.98272, 65.37194, 63.98095, 64.50792,
    65.2442, 67.12506, 70.30002, 72.75606, 73.59404, 71.77447, 58.87996,
    50.49597, 46.43343, 44.96567, 42.87902, 42.17845, 41.8655, 41.28796,
    41.03253, 40.93579,
  66.78082, 65.18594, 63.98185, 63.3516, 63.9224, 64.3358, 64.76099,
    65.08665, 65.39229, 66.10801, 66.16193, 64.82905, 64.73177, 64.9024,
    65.64442, 67.45114, 70.4074, 72.60136, 72.76684, 71.07034, 63.17,
    53.98368, 47.37136, 45.46001, 43.6915, 42.35124, 41.77583, 41.30621,
    41.0199, 40.94283,
  66.09475, 64.77862, 63.47224, 62.85891, 63.31776, 63.6233, 63.98848,
    64.2931, 64.66759, 65.12526, 64.4968, 63.44986, 63.54214, 63.62812,
    64.24072, 65.73656, 66.96481, 64.00092, 63.33956, 62.02201, 59.85451,
    57.35133, 51.89987, 47.63654, 44.76715, 42.96593, 41.72073, 41.28542,
    41.00904, 40.94234,
  66.50497, 64.42728, 63.12521, 62.2534, 62.4583, 62.42037, 62.65624,
    62.75879, 63.25655, 63.29378, 62.13254, 61.42009, 61.41191, 61.50095,
    62.39749, 64.34003, 60.42959, 57.66536, 56.48801, 55.30126, 55.91232,
    56.59196, 54.78149, 53.28956, 48.37837, 43.90903, 41.89149, 41.53706,
    41.05124, 40.93617,
  66.32993, 64.43108, 62.80528, 61.8106, 62.15034, 62.16192, 61.81633,
    61.39933, 61.60258, 61.30322, 60.2831, 60.12751, 60.19834, 60.6451,
    61.75824, 62.7648, 59.4572, 55.31369, 53.32784, 52.50812, 53.15969,
    53.91307, 51.78644, 51.9546, 51.32779, 46.5301, 42.85038, 42.56021,
    41.74941, 41.04103,
  68.12572, 66.31782, 65.07619, 64.31985, 64.33544, 64.0612, 64.11486,
    64.23221, 64.52245, 63.66317, 62.83115, 63.18616, 63.5463, 64.04043,
    64.79728, 66.26385, 62.64342, 58.41014, 54.63305, 53.40745, 53.63074,
    53.17041, 51.22096, 50.04548, 50.10257, 49.81281, 46.28366, 43.24012,
    42.4099, 41.3903,
  70.15354, 70.10133, 67.45108, 66.31746, 66.52669, 66.46342, 66.31851,
    66.61824, 67.37964, 66.71323, 65.48454, 65.87594, 66.33524, 66.65346,
    67.229, 67.74437, 63.08503, 59.57539, 56.09285, 53.28778, 52.813,
    52.21872, 50.59335, 49.2044, 48.16319, 49.01652, 48.82914, 45.76401,
    44.03421, 42.48972,
  72.975, 73.40456, 71.29266, 69.71402, 69.27484, 68.82824, 69.24228,
    69.77811, 69.19867, 67.96106, 67.23884, 67.43973, 67.84923, 67.89666,
    68.19302, 65.61899, 61.89997, 59.19418, 56.56032, 53.91507, 53.56766,
    53.11509, 50.704, 48.737, 48.21773, 48.36829, 49.26517, 47.43676,
    43.83408, 42.26466,
  73.6319, 73.71893, 71.60459, 70.17113, 70.03647, 69.50576, 69.86185,
    69.96062, 68.99562, 68.13689, 67.86094, 67.8933, 67.94197, 67.87904,
    68.47653, 66.23583, 62.70018, 60.80901, 59.09296, 57.67951, 58.71107,
    60.37535, 59.10823, 55.45953, 52.957, 52.0693, 52.6888, 51.22343,
    44.71896, 41.2219,
  73.76112, 73.48267, 71.93124, 71.31255, 71.70979, 71.29832, 70.72794,
    70.02378, 69.05788, 68.87469, 68.73168, 68.8446, 68.87319, 68.82502,
    69.6433, 71.06985, 67.79103, 65.80883, 65.09946, 64.73326, 64.57913,
    62.6923, 58.79651, 56.08714, 54.2779, 53.50238, 52.70963, 54.08494,
    51.12204, 43.35062,
  69.61997, 69.47681, 70.37289, 70.9389, 71.28996, 71.49121, 70.37875,
    68.40654, 67.55131, 67.45108, 67.11496, 66.75332, 66.43386, 66.74286,
    67.97459, 69.73843, 71.19322, 68.42798, 64.41025, 60.25499, 58.27009,
    55.83323, 53.18828, 51.37658, 50.91959, 50.68311, 49.90922, 48.25533,
    47.67427, 44.56963,
  68.45902, 68.42404, 68.66412, 68.58118, 69.05273, 69.91461, 69.62648,
    67.57796, 66.23898, 66.41431, 66.49765, 66.26263, 65.80167, 65.55295,
    66.11168, 67.41872, 64.03311, 57.88612, 55.12489, 52.5698, 50.31869,
    49.28725, 48.39901, 47.62262, 47.15845, 47.15293, 46.6476, 44.9608,
    42.89362, 41.25169,
  26.81858, 26.96123, 27.09664, 27.23097, 27.29139, 27.36932, 27.48856,
    27.63479, 27.83736, 28.08009, 29.02612, 29.20966, 27.87806, 28.01195,
    28.09655, 27.61641, 27.50775, 27.73699, 28.04287, 28.95375, 29.55046,
    29.08327, 29.36086, 30.32584, 31.06218, 30.90799, 33.55936, 35.05379,
    29.25348, 27.1177,
  30.09593, 30.45781, 30.28489, 30.81108, 30.75032, 30.70793, 31.00037,
    31.27938, 31.57276, 31.89536, 32.36737, 33.03642, 33.49576, 32.38597,
    31.38571, 31.19128, 30.23927, 30.43473, 31.30242, 32.2392, 32.49687,
    32.39267, 32.8939, 34.25995, 39.09283, 40.42093, 34.59277, 36.92729,
    29.96526, 27.86808,
  34.40946, 34.83319, 35.0463, 35.41734, 35.71731, 36.05552, 36.39053,
    36.75898, 37.14008, 37.48204, 37.88999, 38.48862, 38.72123, 38.82559,
    38.17576, 36.02077, 35.26241, 35.6307, 35.96949, 36.98465, 38.81599,
    40.85844, 41.78031, 40.92949, 44.55114, 46.71912, 37.88363, 35.87779,
    29.95355, 28.56838,
  41.11346, 41.82622, 42.45924, 43.22145, 43.9588, 44.9928, 45.45911,
    45.51352, 45.88158, 46.42326, 46.80263, 47.2875, 46.81305, 45.18891,
    44.78223, 44.13805, 41.66969, 39.4229, 39.93027, 40.99038, 43.62687,
    44.35018, 41.96494, 46.98419, 49.25525, 41.77727, 40.55488, 34.65409,
    30.08171, 27.68279,
  48.72808, 48.98353, 49.61207, 50.39702, 50.92197, 51.31638, 51.67173,
    51.86508, 52.59821, 53.17609, 52.96203, 52.92486, 52.28259, 51.15567,
    49.20494, 46.99548, 44.11864, 41.36859, 41.1088, 46.42561, 48.53483,
    39.67931, 39.59551, 41.103, 42.91891, 41.88354, 37.92321, 37.78592,
    36.96403, 30.21716,
  53.89244, 54.81176, 55.7319, 57.0313, 56.96195, 56.72715, 57.59186,
    58.13051, 58.19827, 58.89392, 59.74572, 61.90732, 63.59602, 61.14715,
    57.67881, 61.55659, 61.4081, 54.16825, 43.32464, 43.82447, 41.25514,
    37.69576, 38.55646, 39.73856, 41.87766, 40.4287, 44.08278, 56.86537,
    51.25774, 28.7984,
  59.57794, 61.18095, 62.54366, 64.2092, 64.80486, 65.37313, 66.96764,
    67.03385, 66.48677, 66.05901, 65.72319, 64.38371, 60.50578, 58.2802,
    60.86811, 61.60436, 54.94658, 44.73816, 40.69296, 39.96028, 38.38593,
    37.49253, 38.2211, 40.46434, 41.01519, 37.16093, 46.70934, 57.39965,
    47.37852, 26.73644,
  65.39648, 66.24818, 66.7449, 67.11742, 66.86554, 66.78174, 67.1628,
    66.33263, 62.25867, 60.74598, 58.68908, 56.24707, 53.6419, 51.55013,
    49.37809, 46.69331, 43.59084, 41.27666, 38.16341, 37.43732, 36.66579,
    36.61094, 38.17643, 39.88447, 38.69837, 36.47145, 47.68378, 53.25855,
    33.61459, 27.47932,
  65.97851, 66.75045, 67.13731, 67.24141, 66.90307, 66.82083, 63.12323,
    60.39624, 59.97886, 59.17525, 57.94894, 56.65115, 55.22404, 56.9635,
    56.20391, 47.12872, 43.9254, 44.16106, 43.28053, 40.21113, 38.24571,
    40.68038, 45.14444, 45.11189, 40.02806, 40.47757, 43.41081, 39.66529,
    29.53995, 27.2278,
  67.68851, 68.73865, 69.18183, 69.64917, 69.14781, 67.54589, 61.48865,
    62.73664, 63.18712, 64.68018, 66.52682, 68.01014, 67.19626, 62.30786,
    55.21638, 52.87189, 51.32185, 49.6827, 47.15698, 45.84799, 46.26883,
    45.66043, 44.73823, 40.60091, 48.09031, 59.09492, 47.25092, 30.48525,
    27.43223, 26.22348,
  70.43922, 70.96777, 71.73836, 71.60087, 71.64332, 71.44936, 70.81054,
    70.88013, 71.17222, 72.8241, 73.84196, 67.87715, 61.58975, 58.02203,
    54.28156, 51.49669, 49.85683, 48.00084, 45.91393, 44.68889, 46.18083,
    43.87588, 38.33458, 34.65524, 36.34915, 37.55548, 31.64682, 27.11463,
    26.6907, 26.13038,
  75.61572, 72.89684, 76.23443, 77.84261, 77.92952, 76.77583, 75.79886,
    72.74055, 69.55617, 69.86108, 69.03256, 64.28885, 64.69675, 61.99364,
    52.77649, 49.32872, 45.22469, 43.11887, 41.24939, 40.4894, 41.54953,
    39.07818, 33.0371, 37.50396, 40.24387, 29.87246, 26.76936, 27.19306,
    26.94658, 26.38433,
  81.65659, 82.69457, 85.19209, 86.14168, 85.30822, 81.84705, 74.59955,
    70.06162, 70.31287, 68.55503, 68.47044, 67.48137, 66.90067, 65.55883,
    54.90189, 46.8913, 43.48825, 41.24245, 39.55446, 40.7649, 40.67127,
    36.12005, 32.53125, 35.87972, 37.71092, 28.79633, 27.22936, 27.38796,
    27.46673, 26.7517,
  79.07896, 81.0829, 80.53059, 78.60137, 76.58255, 75.13297, 74.63564,
    74.79227, 72.47128, 71.30825, 72.13886, 70.84531, 71.4093, 69.96759,
    65.24248, 56.85408, 44.32632, 45.23989, 45.37543, 44.43204, 38.97727,
    37.97125, 41.05722, 32.47123, 29.08225, 28.10512, 27.27523, 26.90335,
    27.12275, 26.73867,
  71.50415, 71.66714, 71.0285, 70.17523, 69.49172, 71.27418, 76.54415,
    76.95132, 73.86124, 72.98296, 71.83292, 69.84638, 67.87189, 66.86583,
    64.44888, 51.75903, 48.78473, 46.14266, 46.49826, 47.86633, 44.04595,
    36.9474, 31.21941, 29.06103, 28.13947, 28.00193, 27.30385, 26.81121,
    26.63343, 26.37919,
  68.70476, 69.42941, 69.88976, 70.0079, 70.07573, 70.96093, 71.92096,
    71.58324, 70.6347, 69.60679, 69.08442, 67.76618, 64.97665, 62.43072,
    55.01227, 48.65845, 45.86002, 41.70689, 40.32385, 38.86021, 32.81059,
    30.95822, 28.95009, 28.44574, 28.2788, 27.80656, 27.22977, 26.82372,
    26.55449, 26.31511,
  68.31284, 69.01104, 69.28854, 69.53348, 69.92825, 69.54161, 69.61034,
    70.0533, 69.53677, 68.83018, 67.44334, 66.92191, 66.59997, 58.9336,
    50.9664, 45.50988, 41.20866, 37.94948, 38.86488, 37.73418, 30.11516,
    30.30939, 29.35368, 28.49417, 27.9594, 27.80279, 27.17051, 26.54533,
    26.43051, 26.2971,
  67.47265, 68.51352, 68.5075, 68.71149, 68.57036, 68.46632, 68.22188,
    68.35365, 68.61434, 66.68121, 66.41897, 66.9348, 62.08033, 56.59508,
    52.45326, 44.62421, 37.75213, 34.60372, 37.11391, 35.97324, 30.21747,
    30.08779, 29.20966, 28.47854, 27.47946, 27.30984, 27.00554, 26.35962,
    26.25627, 26.1802,
  68.78474, 69.07384, 68.23523, 67.16896, 66.16414, 64.97765, 64.3794,
    64.14539, 62.82333, 61.50089, 62.33748, 59.45415, 51.95474, 48.83003,
    45.40559, 41.77336, 41.07746, 41.79965, 44.19407, 43.23996, 36.82344,
    31.65504, 28.98168, 28.42663, 27.22753, 26.87761, 26.73364, 26.34828,
    26.20686, 26.16066,
  68.74402, 68.76862, 65.21365, 62.22202, 61.22801, 60.42493, 59.79474,
    59.17179, 58.63075, 60.09261, 59.72099, 53.9343, 50.16441, 46.95875,
    43.53756, 40.89692, 41.0291, 42.30687, 43.03771, 42.90382, 39.42422,
    33.68959, 29.25283, 28.53173, 27.63601, 26.96429, 26.64414, 26.35762,
    26.20945, 26.15782,
  67.21472, 65.0174, 61.69275, 59.17048, 58.12194, 57.53259, 57.0743,
    56.76627, 57.18993, 58.67158, 56.56589, 52.05708, 50.40496, 46.99912,
    42.74678, 39.10238, 37.67966, 37.01288, 36.99374, 36.32308, 35.01138,
    33.89855, 31.53746, 29.54461, 28.21119, 27.32225, 26.65987, 26.37589,
    26.21877, 26.16611,
  66.58498, 63.27588, 60.44937, 58.55939, 57.63496, 56.57908, 56.38714,
    56.03299, 57.35699, 57.76367, 54.08097, 50.70657, 48.15566, 43.61266,
    38.96301, 35.87897, 34.10682, 33.17754, 32.79094, 32.02232, 33.34516,
    34.3356, 32.28042, 32.55312, 30.29205, 27.88296, 26.76032, 26.54646,
    26.25512, 26.17019,
  65.50294, 63.29827, 60.23104, 58.55513, 58.77562, 58.60491, 57.59257,
    55.97638, 55.84299, 54.33595, 50.39709, 48.00194, 44.76437, 40.36404,
    36.06157, 34.14397, 33.28946, 31.8858, 31.21004, 30.75145, 32.0686,
    32.82875, 30.35022, 31.42952, 31.69781, 29.23643, 27.22745, 27.18682,
    26.72691, 26.23576,
  65.36948, 63.70938, 62.00314, 61.10744, 60.37991, 59.13981, 58.57649,
    57.51128, 57.02138, 53.40294, 48.94392, 47.51194, 44.62047, 40.82067,
    37.04934, 34.86572, 34.17244, 33.04087, 31.46532, 30.8297, 30.93045,
    30.83057, 30.04435, 29.86786, 30.52484, 30.91431, 29.22377, 27.57336,
    27.10062, 26.4403,
  64.5281, 64.37349, 61.05167, 59.53059, 59.19082, 58.30455, 56.82667,
    55.88298, 56.53518, 53.6618, 49.00227, 48.0218, 45.38719, 41.44063,
    37.76669, 35.8435, 34.52962, 33.85835, 32.63466, 31.13019, 31.02207,
    31.10415, 30.64943, 29.83313, 29.20916, 30.35222, 30.5598, 28.77538,
    27.99695, 27.05145,
  65.19312, 66.37254, 64.16448, 61.27401, 59.34223, 57.97561, 58.28113,
    58.59511, 56.28126, 52.8414, 50.53462, 49.2433, 46.59073, 41.80448,
    37.30156, 35.19439, 34.27227, 33.88387, 33.02703, 31.53407, 31.48968,
    31.56377, 30.36588, 29.40123, 29.3118, 29.74464, 30.7695, 29.86166,
    27.96213, 26.95522,
  66.14391, 66.32213, 62.8807, 60.60857, 59.44567, 57.95842, 58.49062,
    57.88869, 54.48008, 51.90062, 51.03011, 49.40723, 45.92616, 40.87154,
    36.85049, 34.65131, 33.6551, 33.46462, 32.82537, 31.7674, 32.3344,
    33.86024, 33.99456, 32.52725, 31.65594, 31.57721, 32.64506, 32.17747,
    28.35789, 26.31341,
  65.50496, 64.328, 61.81982, 60.91639, 60.49171, 59.132, 58.32137, 55.9353,
    52.12085, 51.19619, 50.10408, 48.25788, 44.72483, 40.12278, 37.04441,
    35.25867, 34.23334, 34.21163, 34.5787, 34.89366, 35.64746, 35.64706,
    34.33089, 33.12879, 32.43025, 32.34169, 32.23186, 33.60717, 32.01582,
    27.46202,
  63.42176, 61.81139, 61.68802, 61.90351, 61.60935, 61.58212, 58.79121,
    53.78694, 51.23586, 50.84445, 49.24392, 46.96136, 43.76599, 40.57075,
    38.63171, 37.63847, 37.4565, 37.71544, 36.58947, 34.81117, 34.25563,
    33.34316, 32.06312, 31.17082, 31.10404, 31.29351, 31.07574, 30.32725,
    30.35902, 28.2778,
  61.34309, 60.88758, 60.11182, 58.79996, 58.32506, 59.88823, 59.62721,
    54.47438, 51.38613, 52.00374, 51.87033, 50.47366, 47.42833, 43.99054,
    41.20956, 39.22632, 37.23327, 35.03141, 33.80312, 32.39083, 31.22781,
    30.66666, 30.21684, 29.78933, 29.57668, 29.75993, 29.58484, 28.64334,
    27.52028, 26.43973,
  25.23559, 25.29886, 25.35098, 25.41047, 25.40232, 25.39989, 25.43293,
    25.47901, 25.5797, 25.70742, 26.49718, 26.63404, 25.64816, 25.79305,
    25.93436, 25.62882, 25.56185, 25.6579, 25.75676, 26.35664, 26.67945,
    26.22576, 26.29139, 26.96297, 27.49339, 27.29288, 29.64516, 31.04271,
    27.30235, 25.87831,
  25.91297, 26.01376, 25.8123, 26.11972, 25.94504, 25.80352, 25.9124,
    26.00504, 26.13689, 26.33091, 26.68272, 27.26743, 27.68447, 26.98904,
    26.63113, 26.79157, 26.32285, 26.49671, 27.08152, 27.64477, 27.71543,
    27.46168, 27.83261, 28.7058, 33.19743, 34.53774, 30.21379, 32.47888,
    27.9346, 26.36214,
  25.99415, 26.04063, 26.04016, 26.11137, 26.13174, 26.18427, 26.27741,
    26.40209, 26.55958, 26.71001, 26.88869, 27.3642, 27.75127, 28.34687,
    28.66528, 27.97871, 28.07332, 28.66587, 28.96652, 29.54095, 30.76721,
    32.29509, 33.40318, 32.81976, 37.46914, 40.27238, 32.48753, 31.93751,
    27.87679, 26.90632,
  26.52135, 26.63935, 26.94499, 27.26078, 27.62983, 28.24348, 28.45527,
    28.31548, 28.47787, 28.86742, 29.06402, 29.52096, 29.60653, 29.39198,
    30.64204, 31.87906, 31.3723, 30.55979, 31.20301, 31.99951, 34.28715,
    35.39318, 33.83791, 38.72375, 41.03412, 35.19784, 34.70893, 31.16321,
    28.00548, 26.31097,
  28.12151, 28.06063, 28.55032, 29.09132, 29.50096, 29.78768, 30.00858,
    30.08451, 30.71081, 31.1368, 30.95341, 31.15697, 31.40099, 31.95915,
    32.74381, 33.48035, 32.96077, 32.34866, 32.69091, 37.62735, 39.33421,
    32.72268, 32.61508, 34.03049, 35.69972, 34.75891, 32.21971, 32.20236,
    32.39452, 28.06281,
  29.5893, 30.10749, 31.03369, 32.12597, 32.07037, 31.73764, 32.25457,
    32.52371, 32.5559, 33.0948, 33.74119, 35.90503, 38.18991, 38.34986,
    37.47415, 46.41923, 56.10527, 43.48093, 35.26313, 36.3376, 34.45414,
    31.34241, 31.83137, 32.60518, 34.6655, 33.58867, 37.3164, 51.99535,
    45.0015, 27.04016,
  31.77586, 32.6913, 33.86348, 35.22928, 35.74375, 36.13378, 37.72704,
    39.81636, 40.37757, 40.38564, 40.92007, 40.10529, 38.36508, 38.00582,
    43.60182, 51.42223, 46.29274, 37.22898, 34.21357, 33.54762, 32.15923,
    31.35824, 31.82025, 33.67847, 34.6652, 31.57441, 41.82744, 58.68124,
    43.17429, 25.56356,
  35.07911, 36.471, 38.13058, 39.8377, 40.24378, 42.09949, 44.08064,
    41.82352, 39.8113, 39.44001, 38.47253, 36.85177, 35.37704, 35.03858,
    36.11982, 37.04045, 35.87751, 34.48301, 32.48141, 31.88644, 31.19714,
    30.97769, 32.13278, 33.59699, 33.1045, 30.94365, 43.2193, 48.92749,
    31.20079, 26.5091,
  40.695, 41.71913, 42.9997, 43.24555, 42.94152, 43.515, 41.411, 39.44414,
    39.13857, 38.54247, 37.34441, 36.06263, 35.32433, 38.503, 40.17216,
    35.68337, 35.02078, 36.16308, 35.76927, 33.24653, 31.47489, 33.0437,
    36.6502, 36.70811, 33.07853, 33.49102, 37.67981, 36.1049, 28.78722,
    26.41889,
  46.49619, 48.45172, 48.98621, 49.40482, 47.58758, 42.89152, 38.0373,
    38.12098, 37.9568, 38.26568, 39.62844, 42.82227, 43.14187, 40.98116,
    38.3249, 38.34861, 38.72758, 38.39452, 36.99316, 36.59659, 37.02941,
    37.33816, 37.47793, 34.82766, 41.95702, 53.18478, 42.11023, 29.21808,
    26.776, 25.3811,
  60.35005, 58.89776, 59.16837, 53.81363, 51.33973, 48.25713, 44.52598,
    46.40535, 47.7064, 57.22525, 64.43916, 43.25296, 37.80307, 36.88394,
    36.16667, 36.94777, 38.55033, 37.97188, 36.59326, 36.245, 38.68175,
    37.80779, 33.75946, 30.96783, 34.06158, 36.87875, 31.10314, 26.30469,
    25.78146, 25.24472,
  64.24354, 58.6478, 61.32042, 62.26638, 63.10958, 62.67632, 62.79326,
    56.82444, 46.64494, 49.69481, 48.85641, 36.9211, 38.92793, 39.9925,
    36.80093, 37.03616, 35.9756, 35.29848, 34.23138, 34.29922, 36.69642,
    35.07039, 29.90759, 34.22099, 36.29495, 28.38553, 25.78531, 26.17568,
    26.04951, 25.49347,
  68.04454, 66.5276, 71.13829, 72.23259, 73.16954, 70.60023, 63.28673,
    49.89808, 49.43892, 45.3309, 43.81209, 38.94484, 42.96375, 44.39815,
    37.71764, 36.72692, 36.12835, 34.7405, 33.33846, 35.3635, 36.51201,
    32.62252, 29.32798, 34.21886, 35.74001, 27.57701, 26.11444, 26.34562,
    26.60029, 25.8206,
  70.22227, 74.51286, 73.04203, 70.79436, 68.25928, 64.98807, 61.73397,
    61.4054, 60.94433, 61.11634, 64.69169, 68.90524, 69.97291, 66.8138,
    56.79446, 44.02497, 35.99548, 37.56384, 38.60647, 39.14231, 35.40593,
    34.50742, 36.47175, 30.75246, 28.19953, 26.89003, 26.13612, 25.85579,
    26.25879, 25.78802,
  64.69869, 63.86552, 62.396, 60.7028, 59.04537, 59.67278, 64.0158, 64.40479,
    62.21201, 61.97963, 64.29801, 57.94965, 45.9845, 51.42213, 55.22162,
    40.01011, 39.90892, 39.31732, 42.24988, 43.92529, 39.18198, 34.24642,
    29.83502, 27.49142, 26.71584, 26.92266, 26.2593, 25.78518, 25.71313,
    25.46202,
  58.14527, 55.83107, 54.81107, 53.90361, 54.6706, 58.63171, 59.74867,
    59.84681, 57.1414, 53.18284, 48.54883, 42.44258, 39.77463, 42.35103,
    41.21107, 38.80611, 39.52148, 37.28059, 37.88494, 37.40328, 31.40839,
    28.95529, 27.07694, 26.84445, 27.04933, 26.79636, 26.29621, 25.86412,
    25.63443, 25.38159,
  53.97196, 51.99057, 50.97102, 50.58099, 50.82935, 50.06347, 48.97724,
    47.98109, 45.95378, 43.57924, 39.96275, 41.24184, 45.34472, 42.04887,
    38.9316, 37.9894, 36.46622, 34.27928, 36.50149, 35.46207, 27.90629,
    28.14704, 27.64739, 26.96943, 26.71722, 26.79677, 26.24282, 25.604,
    25.51023, 25.36499,
  49.68726, 48.70524, 47.28303, 46.47308, 45.27184, 44.52924, 44.01923,
    43.48161, 42.43301, 40.39659, 40.89085, 43.77141, 42.75164, 41.84692,
    42.61214, 38.92356, 33.82869, 31.25525, 34.66861, 33.75619, 28.16731,
    28.34518, 27.91854, 27.23498, 26.30535, 26.34557, 26.04464, 25.43498,
    25.33775, 25.27205,
  48.23919, 46.58208, 43.80545, 41.86169, 41.03619, 40.17808, 39.80375,
    39.80162, 38.89661, 38.21254, 40.43943, 39.73807, 35.13665, 35.55362,
    36.02065, 34.85943, 34.82356, 35.53856, 38.84068, 38.41389, 32.83503,
    29.53221, 28.05799, 27.35116, 26.16588, 25.93578, 25.7951, 25.42814,
    25.30665, 25.25477,
  45.33933, 43.47312, 40.98219, 38.9228, 38.26988, 37.75578, 37.37681,
    36.98162, 36.61266, 38.64384, 39.02723, 34.36323, 32.38092, 32.59202,
    32.52859, 32.01247, 33.40253, 35.4703, 37.50665, 38.66221, 36.02221,
    31.47865, 28.27654, 27.43822, 26.55454, 25.98057, 25.71453, 25.43909,
    25.30282, 25.25129,
  42.45139, 41.41865, 39.09678, 37.19481, 36.37333, 35.88454, 35.34447,
    34.83081, 35.18777, 37.06223, 35.00709, 31.22295, 32.04184, 32.75133,
    32.49105, 31.56792, 31.55717, 31.81062, 32.89042, 33.27698, 32.70664,
    32.04674, 30.24183, 28.26878, 27.03142, 26.26905, 25.70724, 25.44064,
    25.319, 25.2629,
  41.18305, 39.59943, 37.46523, 36.09776, 35.22342, 34.09775, 33.69868,
    33.31514, 34.93591, 35.78541, 32.57854, 30.79428, 31.728, 31.90474,
    31.44735, 30.84434, 30.10058, 29.62295, 29.62348, 29.25501, 30.82937,
    31.66444, 31.03258, 31.5569, 29.29898, 26.8787, 25.85315, 25.62377,
    25.36165, 25.26359,
  40.08816, 38.23671, 35.87232, 34.57999, 34.94993, 35.11144, 34.564,
    33.72008, 34.84014, 34.2104, 31.07593, 30.56503, 30.85972, 30.8161,
    30.19599, 30.32729, 30.06554, 28.83703, 28.33589, 28.12121, 29.78834,
    30.24034, 28.71729, 30.38268, 30.75744, 28.13801, 26.26352, 26.26794,
    25.78212, 25.3143,
  39.13095, 37.41888, 36.49259, 36.18606, 36.14979, 36.05309, 36.49465,
    36.57694, 37.35495, 34.42282, 30.63728, 30.82483, 31.16507, 31.45353,
    31.1538, 30.89796, 30.97038, 30.03543, 28.62339, 28.28221, 28.7415,
    28.70344, 28.08427, 28.29718, 29.51286, 29.94654, 28.13526, 26.63065,
    26.15269, 25.49432,
  38.81064, 39.08699, 36.75515, 35.98876, 36.40321, 36.38175, 35.8171,
    35.78401, 37.29729, 34.54299, 30.45808, 30.92188, 31.5291, 31.65536,
    31.57428, 31.58506, 31.13219, 30.90035, 29.66864, 28.24055, 28.52018,
    28.83157, 28.6183, 27.863, 27.40176, 28.8656, 29.12903, 27.52987,
    27.04328, 26.01077,
  39.90581, 41.52751, 40.34468, 38.33379, 36.83064, 35.84314, 36.71704,
    37.76207, 36.20533, 33.07649, 31.14283, 31.64728, 32.39745, 31.85583,
    31.01624, 30.94125, 30.76088, 30.7888, 30.01839, 28.5718, 29.05847,
    29.47051, 28.32413, 27.39167, 27.24888, 27.82594, 29.22233, 28.3746,
    26.91467, 25.87764,
  41.0375, 41.83145, 39.0058, 37.13016, 36.19132, 35.21285, 36.56922,
    36.95301, 33.90132, 31.63635, 31.43319, 31.84498, 32.05598, 31.38746,
    30.87902, 30.54041, 30.22937, 30.40612, 29.7461, 28.4996, 29.44157,
    31.38639, 31.62622, 30.06483, 29.18305, 29.24139, 30.76832, 30.4105,
    27.02514, 25.29532,
  40.18396, 39.55474, 37.55371, 36.94849, 37.17363, 36.60962, 36.96473,
    35.35646, 31.83953, 31.2274, 31.06866, 31.39105, 31.44119, 30.98955,
    31.15414, 30.88756, 30.2275, 30.33717, 30.60922, 30.64892, 32.1892,
    32.88992, 31.74464, 30.31661, 29.61774, 29.72653, 29.93505, 31.82538,
    30.222, 26.19271,
  37.58918, 36.30349, 36.67175, 37.75806, 38.58299, 39.5134, 37.69376,
    33.52814, 31.31365, 31.10439, 30.11469, 29.68903, 29.70351, 30.29096,
    31.39408, 31.95003, 32.31303, 33.02089, 32.0209, 30.55737, 30.64785,
    30.08248, 28.88474, 28.15146, 28.23844, 28.71961, 28.82146, 28.53444,
    28.96734, 26.85181,
  36.9508, 36.87803, 36.6022, 36.08508, 36.38112, 38.86174, 39.34819,
    34.43999, 31.42699, 31.94059, 32.28746, 32.71809, 32.99319, 33.6139,
    34.20148, 34.12255, 32.88368, 31.24511, 30.22272, 28.9262, 28.13688,
    27.79487, 27.48912, 27.26177, 27.24501, 27.73352, 27.85123, 27.1626,
    26.39349, 25.5011,
  22.93352, 22.98445, 23.04159, 23.08032, 23.06838, 23.05092, 23.05357,
    23.08599, 23.14063, 23.22974, 24.13223, 24.20782, 23.22772, 23.39261,
    23.5057, 23.19031, 23.10299, 23.15448, 23.18358, 23.77289, 24.05269,
    23.52398, 23.52531, 24.13557, 24.50186, 24.14065, 26.72201, 28.35721,
    25.00513, 23.64108,
  23.45168, 23.49184, 23.2906, 23.57364, 23.36674, 23.20648, 23.27532,
    23.32619, 23.41531, 23.58419, 23.97788, 24.56702, 24.93731, 24.2104,
    23.88792, 23.95704, 23.43961, 23.49938, 24.01872, 24.56389, 24.5283,
    24.03656, 24.15713, 25.04125, 29.26408, 29.81514, 27.4136, 30.4268,
    25.80358, 24.21199,
  23.37545, 23.39534, 23.36053, 23.40763, 23.36185, 23.33989, 23.37013,
    23.44899, 23.55214, 23.61951, 23.74742, 24.19847, 24.53135, 25.10737,
    25.28164, 24.41662, 24.34696, 24.75312, 24.83859, 25.22275, 26.23396,
    27.66374, 28.74734, 28.3794, 33.03483, 35.30275, 29.841, 29.90314,
    25.735, 24.7508,
  23.52577, 23.53248, 23.74386, 23.92914, 24.21912, 24.77152, 24.85296,
    24.58994, 24.62685, 24.89935, 25.05471, 25.46053, 25.31414, 25.01758,
    26.16435, 27.26191, 26.54912, 25.52922, 25.86313, 26.47755, 29.11195,
    30.37517, 29.23349, 33.85428, 35.48209, 31.85858, 32.45891, 29.39672,
    25.88282, 24.10697,
  24.33634, 24.12458, 24.4346, 24.82765, 25.14403, 25.37032, 25.44684,
    25.32218, 25.89022, 26.254, 25.99314, 26.00588, 26.00957, 26.45216,
    27.2566, 27.894, 27.19584, 26.47584, 26.99823, 32.1156, 33.58928,
    28.11009, 27.89163, 29.72454, 31.65962, 31.16731, 29.38645, 29.87931,
    30.54686, 25.89318,
  24.85912, 25.0874, 25.94856, 27.01883, 26.82233, 26.32341, 26.64047,
    26.55556, 26.2408, 26.42711, 26.63692, 28.79998, 31.19346, 31.29206,
    30.80927, 38.10434, 45.12659, 36.22355, 30.09979, 32.01344, 30.10862,
    26.57285, 27.04474, 27.95517, 30.68868, 30.03951, 32.89792, 45.59071,
    40.51664, 25.07257,
  25.80305, 26.2905, 27.21464, 28.29778, 28.46467, 28.38588, 29.62208,
    31.44739, 31.75767, 31.77108, 32.60044, 32.2471, 31.01159, 31.13619,
    36.83811, 43.81801, 40.2005, 32.42113, 29.47528, 29.01431, 27.46945,
    26.47789, 27.07701, 29.57693, 30.96691, 28.20314, 38.57819, 53.94963,
    39.9836, 23.56411,
  27.06038, 27.78266, 29.05627, 30.39671, 30.59743, 32.84089, 35.35328,
    33.38415, 31.76192, 31.79686, 31.46816, 30.22277, 29.01927, 29.06715,
    31.08773, 32.46618, 31.15588, 29.63672, 27.74795, 27.26255, 26.61408,
    26.42928, 27.82939, 30.07288, 29.61168, 27.98474, 40.74178, 45.62642,
    29.77303, 23.93418,
  30.30412, 31.06902, 32.65257, 33.18619, 33.74263, 35.47711, 34.12674,
    32.3903, 32.31895, 32.01344, 30.90883, 29.54228, 28.68925, 32.34092,
    34.45386, 30.39131, 29.83338, 31.3636, 31.30238, 28.7595, 26.70167,
    28.32447, 32.64871, 33.11113, 29.43975, 29.99575, 36.3973, 34.52351,
    26.02654, 23.90465,
  35.36739, 37.68879, 39.80748, 41.64676, 40.91299, 36.29618, 31.71303,
    31.54099, 31.01911, 30.49927, 31.54617, 35.12469, 36.2452, 34.80522,
    32.75863, 32.71136, 33.26992, 33.71099, 32.25966, 30.61955, 30.77944,
    31.51158, 32.32955, 30.27372, 35.99954, 46.16595, 38.32164, 26.98283,
    24.37452, 23.16528,
  49.63622, 52.53711, 48.48712, 42.60461, 40.77365, 39.19947, 35.31865,
    37.0635, 38.58102, 47.00232, 51.71681, 36.06139, 31.52843, 30.63654,
    29.92336, 30.81477, 31.97854, 31.801, 30.54449, 30.43421, 33.10952,
    32.77457, 29.44794, 27.17834, 31.01369, 34.70921, 28.91159, 23.94282,
    23.52104, 23.03105,
  62.79528, 51.95219, 55.96439, 58.40779, 56.29534, 48.04395, 49.7719,
    46.07881, 38.82222, 42.85601, 42.38826, 29.83739, 30.94993, 31.90055,
    29.98426, 30.35737, 29.74452, 29.54433, 28.92649, 29.43825, 32.32059,
    31.0571, 26.70263, 30.73054, 32.46283, 25.93039, 23.55703, 23.87198,
    23.72272, 23.19675,
  72.18882, 71.14641, 91.83627, 96.71848, 94.29305, 81.05227, 60.88992,
    41.22393, 39.90913, 37.20668, 34.59498, 29.34707, 33.88605, 36.2017,
    31.55429, 30.29103, 30.40197, 29.69903, 28.63703, 30.8074, 32.33199,
    29.14971, 26.17296, 31.64352, 32.77182, 25.21543, 23.77549, 24.00646,
    24.23428, 23.46442,
  80.0319, 97.37112, 99.07665, 95.50202, 80.03717, 69.96083, 66.99718,
    62.39808, 52.27241, 48.11365, 55.58741, 54.31212, 56.48185, 54.36526,
    47.08302, 36.96058, 30.91894, 32.50902, 33.67342, 34.61671, 31.63937,
    30.78783, 32.33094, 28.43422, 26.10911, 24.4857, 23.78792, 23.55705,
    23.97618, 23.4463,
  59.37421, 64.34982, 60.13317, 55.56069, 49.13212, 57.17784, 80.64406,
    78.00769, 68.29162, 68.17274, 65.22614, 50.56398, 40.56471, 45.73235,
    47.22647, 34.34415, 34.69765, 34.77758, 38.20422, 39.14285, 34.5121,
    30.98975, 27.64822, 25.08076, 24.23434, 24.55947, 23.91158, 23.46408,
    23.44235, 23.18432,
  46.01502, 44.1256, 42.6757, 41.06351, 41.38657, 47.36555, 54.42791,
    52.74585, 49.76719, 47.45271, 43.91497, 36.84237, 32.65212, 36.23142,
    35.9229, 33.57642, 35.11526, 33.68582, 35.06501, 34.50547, 28.86337,
    26.34118, 24.3869, 24.22506, 24.60525, 24.44913, 23.9789, 23.54488,
    23.38236, 23.11445,
  41.40653, 39.27633, 38.35857, 38.42818, 39.77996, 40.69705, 41.01922,
    41.02197, 39.78148, 37.69829, 33.71476, 33.95547, 38.27782, 36.06261,
    33.75363, 33.56308, 32.85009, 31.22136, 33.538, 31.99388, 25.17729,
    25.30519, 24.86927, 24.29823, 24.26163, 24.39719, 23.87188, 23.32623,
    23.28928, 23.10768,
  37.42871, 37.08439, 36.84232, 37.40977, 37.49418, 37.83889, 37.65713,
    37.27889, 36.60371, 33.71413, 33.81667, 37.1391, 37.33067, 36.83207,
    37.83958, 35.06083, 30.69403, 28.47768, 31.88307, 30.41594, 25.36153,
    25.61873, 25.28134, 24.59112, 23.85158, 24.01655, 23.68272, 23.15687,
    23.11244, 23.02665,
  38.17037, 38.158, 36.62651, 35.65226, 35.30064, 34.65952, 34.19262,
    33.92101, 32.85322, 31.7423, 34.5341, 34.9144, 31.00794, 31.78294,
    32.41995, 31.27621, 31.08974, 31.76591, 35.18396, 34.39222, 29.36697,
    26.70111, 25.52703, 24.80473, 23.77047, 23.633, 23.49289, 23.1504,
    23.06602, 23.00668,
  38.51657, 37.88909, 35.74458, 33.75127, 33.18139, 32.66098, 32.2549,
    31.83523, 31.44283, 33.57628, 34.42708, 30.39125, 28.32812, 28.62071,
    28.40045, 27.87664, 29.45825, 31.81347, 34.33897, 35.35852, 32.61765,
    28.48004, 25.70702, 24.90322, 24.12915, 23.64788, 23.43112, 23.17629,
    23.07561, 23.01145,
  37.12148, 36.22799, 34.19071, 32.46643, 31.81981, 31.55707, 31.26918,
    30.8721, 31.19646, 33.1274, 30.98455, 27.05188, 27.59508, 28.21305,
    27.92152, 27.28452, 27.66357, 28.42542, 29.97481, 30.41774, 29.76847,
    29.05752, 27.41181, 25.61717, 24.56219, 23.89865, 23.42524, 23.18259,
    23.09983, 23.01669,
  36.7218, 34.737, 33.10209, 32.01017, 31.42797, 30.72813, 30.3805, 29.86447,
    31.09344, 31.4513, 27.92537, 26.10056, 27.13998, 27.51419, 27.30961,
    27.00388, 26.58532, 26.45122, 26.68127, 26.48162, 27.58015, 28.17402,
    28.3646, 28.65069, 26.61662, 24.39985, 23.56371, 23.34067, 23.15242,
    23.03255,
  35.57441, 34.1261, 32.17284, 31.10871, 31.41172, 31.482, 30.83191,
    29.76598, 30.58439, 29.54056, 26.3953, 26.03098, 26.65787, 26.90857,
    26.56624, 26.87292, 26.64661, 25.66467, 25.34945, 25.31935, 26.55711,
    26.75864, 26.28126, 27.94267, 28.06124, 25.40574, 23.87904, 23.87936,
    23.49035, 23.07933,
  34.51623, 33.36163, 32.53188, 32.16082, 32.04132, 31.95482, 32.18947,
    32.0048, 32.59139, 29.66688, 26.2757, 26.63427, 27.24096, 27.7794,
    27.60645, 27.50303, 27.66427, 26.80387, 25.6268, 25.50382, 25.90404,
    25.76821, 25.40683, 25.81384, 27.0417, 27.11591, 25.44273, 24.23623,
    23.85071, 23.20748,
  33.8838, 34.05603, 32.16933, 31.6269, 32.11273, 32.11493, 31.59207,
    31.67175, 33.16465, 30.14633, 26.35964, 26.93705, 27.72297, 28.02916,
    28.05593, 28.08119, 27.85196, 27.65888, 26.47655, 25.35843, 25.7009,
    25.90015, 25.70408, 25.04108, 24.82573, 26.23826, 26.38564, 25.00838,
    24.69127, 23.58221,
  34.00755, 35.75011, 35.06307, 33.42138, 32.41909, 31.7, 32.5601, 33.5808,
    32.28426, 28.99993, 26.93699, 27.5793, 28.50301, 28.12273, 27.48524,
    27.47829, 27.38483, 27.54701, 26.77251, 25.60135, 26.19839, 26.47221,
    25.36348, 24.57023, 24.51706, 25.14332, 26.64769, 25.72178, 24.53825,
    23.44765,
  35.21215, 36.57603, 34.28155, 32.63477, 31.98118, 31.32021, 32.79486,
    33.21899, 30.10742, 27.6005, 27.21184, 27.79298, 28.2033, 27.75796,
    27.34501, 27.10469, 26.94531, 27.20221, 26.56968, 25.53496, 26.55231,
    28.19346, 28.04461, 26.63459, 26.17281, 26.36989, 28.21398, 27.66946,
    24.5105, 22.96353,
  34.82806, 34.77897, 33.05038, 32.61808, 33.13114, 32.94101, 33.59698,
    31.72813, 27.95177, 27.06609, 26.90771, 27.41191, 27.69326, 27.49387,
    27.73331, 27.4291, 26.84406, 27.03487, 27.23829, 27.2411, 28.84675,
    29.29321, 28.10544, 26.78761, 26.56903, 26.78214, 27.31848, 29.3259,
    27.41214, 23.7004,
  32.63528, 31.69472, 32.24508, 33.55893, 34.85055, 36.19502, 34.47099,
    30.09641, 27.54831, 27.05552, 26.12402, 25.876, 26.08479, 26.7515,
    27.81124, 28.21966, 28.47544, 29.15539, 28.1998, 27.05813, 27.27119,
    26.74759, 25.61279, 25.039, 25.28901, 25.86898, 26.06145, 26.07269,
    26.65068, 24.26208,
  32.08339, 32.25746, 32.30152, 32.1955, 32.88047, 35.66916, 35.881, 30.6333,
    27.55333, 27.61937, 27.76241, 28.26537, 28.73805, 29.47477, 30.06951,
    30.05628, 28.88267, 27.57858, 26.71957, 25.59691, 24.94815, 24.71867,
    24.49922, 24.3833, 24.47639, 25.11497, 25.27704, 24.65383, 24.08983,
    23.22243,
  15.92872, 15.9615, 16.00493, 16.03635, 16.01329, 16.00263, 16.01044,
    16.01894, 16.06747, 16.11461, 16.86373, 16.89518, 16.12838, 16.30366,
    16.38747, 16.09594, 16.02597, 16.0614, 16.06763, 16.52804, 16.7345,
    16.30591, 16.27842, 16.77105, 17.04583, 16.67798, 18.9272, 20.21866,
    17.64721, 16.53113,
  16.28652, 16.28733, 16.14591, 16.37308, 16.19455, 16.05818, 16.11772,
    16.15856, 16.21573, 16.34617, 16.70477, 17.23446, 17.57673, 16.91971,
    16.6413, 16.63445, 16.20262, 16.22452, 16.60159, 17.00393, 16.96084,
    16.50412, 16.57002, 17.21457, 21.10812, 21.39913, 19.51457, 22.18629,
    18.55387, 17.02842,
  16.20382, 16.20633, 16.17682, 16.21154, 16.15738, 16.12366, 16.14643,
    16.21069, 16.28628, 16.33413, 16.43192, 16.83595, 17.13777, 17.58243,
    17.60922, 16.84343, 16.73926, 16.99048, 17.01251, 17.21846, 17.9355,
    19.09315, 20.10823, 19.6732, 24.25599, 26.21242, 21.94043, 22.37777,
    18.45097, 17.47435,
  16.22412, 16.21648, 16.36632, 16.48359, 16.7091, 17.13428, 17.17794,
    16.94529, 16.98482, 17.24743, 17.31654, 17.61664, 17.42645, 17.18555,
    18.03635, 18.87206, 18.20018, 17.28589, 17.46785, 17.80291, 20.07533,
    21.25958, 20.46373, 24.70575, 26.03833, 23.76054, 24.95039, 22.03798,
    18.46368, 16.91436,
  16.65982, 16.47752, 16.69525, 17.00112, 17.27143, 17.44663, 17.46284,
    17.32772, 17.85988, 18.17007, 17.90381, 17.7706, 17.63022, 17.87554,
    18.53222, 19.05953, 18.27847, 17.67295, 18.09831, 22.66624, 23.86295,
    19.55728, 19.47383, 21.36226, 22.93559, 22.83, 22.02687, 22.44128,
    22.93958, 18.54085,
  16.85821, 16.97693, 17.71483, 18.64279, 18.46153, 17.98698, 18.12667,
    17.93817, 17.63441, 17.72059, 17.69779, 19.44989, 21.36018, 21.44065,
    20.79097, 27.36176, 33.21455, 25.73671, 20.96021, 23.05742, 21.48042,
    18.35668, 18.83731, 19.47183, 21.92951, 21.40112, 24.44901, 36.21332,
    31.86432, 17.92743,
  17.50389, 17.85231, 18.627, 19.49532, 19.48381, 19.14466, 19.94222,
    21.34951, 21.557, 21.53086, 22.3188, 22.07547, 21.13411, 21.20455,
    25.94548, 32.61585, 30.44017, 23.2983, 20.86123, 20.51162, 19.13869,
    18.27427, 18.83902, 21.1441, 22.42668, 19.76137, 29.23238, 43.06755,
    30.9483, 16.56286,
  18.61643, 19.03708, 19.97617, 20.93427, 20.85571, 22.6772, 24.65388,
    22.84178, 21.52687, 21.60231, 21.50971, 20.51821, 19.59893, 19.72437,
    21.94254, 23.56713, 22.35806, 20.82806, 19.39527, 18.9966, 18.45978,
    18.34121, 19.61171, 21.9116, 21.60008, 19.99871, 32.29557, 36.64585,
    22.31407, 16.75999,
  21.42961, 21.83922, 23.06507, 23.34347, 23.83789, 25.45853, 24.37757,
    22.56932, 22.20532, 21.96647, 21.17544, 20.12493, 19.44328, 22.69409,
    24.4388, 21.20813, 21.13, 22.6517, 22.59027, 20.27609, 18.44646,
    19.88416, 23.86347, 24.37349, 21.24104, 21.7723, 28.4567, 26.639,
    18.79304, 16.78504,
  25.6844, 27.39595, 29.15388, 30.50835, 30.41632, 26.99419, 23.25251,
    22.61915, 21.74066, 20.71139, 21.47819, 24.50061, 25.82273, 25.33993,
    23.91462, 23.80252, 24.53877, 25.16112, 23.75798, 22.08655, 22.00087,
    22.83739, 23.91032, 22.40873, 27.33, 36.14332, 29.73215, 19.7178,
    17.27548, 16.15813,
  36.99681, 40.32623, 37.5711, 32.92954, 31.70792, 30.09208, 26.46589,
    27.4754, 28.07592, 34.88198, 37.99918, 25.96793, 22.67465, 22.01393,
    21.32876, 22.29805, 23.51052, 23.39155, 22.10297, 21.88012, 24.22212,
    24.07536, 21.25005, 19.42309, 23.42962, 27.39299, 21.81812, 16.90269,
    16.47459, 16.02232,
  49.54489, 41.19886, 43.18333, 44.57826, 42.7595, 37.33407, 39.46313,
    36.06938, 29.3494, 33.34973, 32.81502, 20.88496, 21.81411, 22.63673,
    21.17003, 21.59039, 21.19412, 20.99706, 20.38519, 20.97611, 23.79978,
    22.75291, 18.99346, 22.40777, 23.83367, 18.50644, 16.43708, 16.78543,
    16.67397, 16.1692,
  56.62111, 53.85459, 69.57092, 75.93508, 74.85446, 65.67192, 50.56668,
    33.72318, 30.41867, 28.48061, 25.50693, 19.43265, 23.88873, 26.2559,
    22.37571, 21.55457, 21.78308, 20.93861, 20.18034, 22.44393, 24.07652,
    21.27918, 18.62257, 23.70483, 24.5405, 17.92421, 16.62886, 16.90445,
    17.13396, 16.40422,
  64.11769, 89.98586, 90.7371, 87.49793, 77.55785, 66.17424, 55.09761,
    49.64048, 40.37782, 35.65347, 41.02378, 39.39643, 41.84538, 41.07967,
    35.32121, 27.03446, 22.14106, 23.4211, 24.63537, 25.86355, 23.44674,
    22.69804, 23.98064, 21.00386, 18.84469, 17.22514, 16.68137, 16.5167,
    16.91775, 16.3847,
  49.19087, 57.62037, 55.96975, 53.31022, 46.92263, 49.36586, 65.38078,
    63.64914, 53.10222, 53.31655, 51.5826, 39.42741, 30.74801, 35.56673,
    36.60577, 25.51551, 25.14984, 25.48839, 28.27671, 29.48261, 26.27584,
    23.27623, 20.5571, 17.93938, 16.91372, 17.25422, 16.75519, 16.38592,
    16.4166, 16.16358,
  38.34093, 38.03181, 37.03839, 35.2729, 34.24873, 38.72813, 45.57944,
    43.5671, 39.84451, 38.36422, 35.29436, 27.68184, 23.39968, 27.10915,
    26.67702, 24.4143, 25.94368, 24.77856, 26.00143, 25.79076, 21.60298,
    19.17951, 17.18665, 17.04968, 17.31132, 17.12777, 16.78028, 16.46123,
    16.34045, 16.09939,
  35.55849, 34.09834, 32.46571, 31.73263, 32.55578, 33.41951, 33.57646,
    33.09991, 31.54785, 29.05952, 24.76885, 24.17167, 27.2579, 25.86042,
    24.54278, 24.58491, 24.22889, 22.79865, 24.32527, 22.95782, 17.82989,
    17.89654, 17.61295, 17.18225, 17.05626, 17.10051, 16.6925, 16.27622,
    16.26364, 16.0884,
  31.72047, 30.81429, 30.03931, 30.57214, 30.97516, 31.54342, 31.49442,
    30.80133, 29.20796, 25.41711, 24.34826, 27.08568, 27.65954, 27.4754,
    28.64657, 26.39547, 22.71602, 20.685, 23.21641, 21.78049, 17.92533,
    18.19709, 18.01878, 17.44594, 16.72915, 16.82869, 16.54635, 16.13588,
    16.10884, 16.02617,
  31.28238, 31.2344, 30.03851, 29.64061, 29.75478, 29.44958, 28.93206,
    27.95077, 25.72231, 23.5537, 25.58326, 26.09034, 23.07477, 23.99984,
    24.66893, 23.45568, 22.97479, 23.32883, 25.67755, 24.68515, 21.08058,
    19.1359, 18.21264, 17.59435, 16.66223, 16.53121, 16.40975, 16.13717,
    16.06656, 16.00231,
  31.88263, 31.82383, 30.17946, 28.7057, 28.46845, 27.97079, 27.23234,
    26.11582, 24.6212, 25.54708, 26.14356, 22.71782, 20.7785, 20.95631,
    20.64908, 20.08897, 21.3953, 23.45925, 25.35333, 26.00309, 24.05889,
    20.70921, 18.31983, 17.64655, 16.95947, 16.55348, 16.36633, 16.15138,
    16.07878, 16.00784,
  31.45429, 31.28673, 29.52332, 27.96117, 27.44198, 27.19874, 26.69729,
    25.7608, 25.19014, 26.18769, 23.84041, 19.90041, 20.06888, 20.32824,
    19.84674, 19.32876, 19.78877, 20.6242, 21.87591, 22.21708, 21.95068,
    21.39928, 19.79278, 18.2028, 17.32239, 16.75576, 16.37263, 16.14905,
    16.08848, 16.01564,
  31.75738, 30.44033, 28.84106, 27.83968, 27.437, 26.93843, 26.63019,
    25.70973, 25.76245, 25.06495, 21.05721, 18.65196, 19.34222, 19.6803,
    19.54094, 19.3274, 19.00817, 18.91383, 19.18845, 19.0341, 20.03417,
    20.30904, 20.08249, 20.39637, 18.92036, 17.11088, 16.47504, 16.26347,
    16.11274, 16.02188,
  31.27835, 30.23812, 28.36417, 27.52816, 28.01069, 28.20253, 27.56985,
    25.95261, 25.47198, 23.22845, 19.33426, 18.38951, 18.92899, 19.25813,
    19.03012, 19.25583, 18.99859, 18.1886, 17.97786, 17.95501, 19.06467,
    18.95974, 18.33566, 20.00154, 20.19498, 17.87825, 16.67841, 16.66706,
    16.36809, 16.05347,
  30.57654, 29.85485, 28.99445, 28.76107, 28.8935, 28.956, 28.83712,
    27.75175, 26.86436, 22.94131, 19.04499, 18.98507, 19.58081, 20.06973,
    19.85293, 19.78704, 19.82984, 19.02148, 18.1616, 18.13223, 18.39182,
    18.15945, 17.82946, 18.27389, 19.37246, 19.46379, 18.05158, 17.00636,
    16.71866, 16.16626,
  30.45525, 31.00151, 29.03075, 28.38687, 28.78261, 28.68758, 27.95773,
    27.32674, 27.45168, 23.3824, 19.21312, 19.30649, 19.92422, 20.28245,
    20.27788, 20.22391, 19.92807, 19.6263, 18.77809, 18.03184, 18.15078,
    18.22664, 18.11734, 17.60654, 17.56595, 18.88281, 18.93371, 17.68837,
    17.53115, 16.49431,
  30.79589, 32.78077, 31.32802, 29.5824, 28.64493, 27.93576, 28.41135,
    28.7702, 26.79434, 22.5384, 19.72269, 19.81662, 20.47268, 20.2468,
    19.75605, 19.7128, 19.47801, 19.45193, 18.9859, 18.18908, 18.46647,
    18.60234, 17.81232, 17.2706, 17.26284, 17.88497, 19.18464, 18.29749,
    17.49697, 16.41885,
  31.62492, 33.33495, 30.81865, 29.00188, 28.25686, 27.57204, 28.80031,
    28.77521, 24.9218, 21.17597, 19.95045, 20.04461, 20.27052, 19.93608,
    19.57717, 19.34921, 19.09367, 19.19543, 18.82998, 18.13652, 18.63482,
    19.79787, 19.71587, 18.88976, 18.75806, 18.88053, 20.62418, 20.06623,
    17.37295, 16.01065,
  31.07352, 31.45624, 29.46598, 28.89731, 29.37358, 29.11042, 29.56614,
    27.30132, 22.79554, 20.5116, 19.59187, 19.63893, 19.76765, 19.73885,
    19.98007, 19.6396, 19.02043, 19.02989, 19.34247, 19.54333, 20.4015,
    20.51948, 19.84137, 19.1082, 19.16627, 19.20459, 19.79125, 21.60276,
    19.79038, 16.57809,
  28.8492, 28.20091, 28.71919, 30.00898, 31.19461, 32.18598, 30.47256,
    25.80233, 22.11988, 20.3885, 18.8459, 18.32731, 18.49924, 18.96709,
    19.71798, 19.99137, 20.08018, 20.58473, 20.08416, 19.45181, 19.56542,
    19.08436, 18.15869, 17.72884, 18.0084, 18.47531, 18.60071, 18.75441,
    19.33593, 17.04006,
  27.92997, 28.22279, 28.49954, 28.66821, 29.19047, 31.54868, 31.18153,
    25.61412, 21.66312, 20.48448, 19.82633, 20.00396, 20.48944, 20.84321,
    21.08133, 21.17618, 20.38071, 19.53984, 19.02454, 18.19116, 17.67065,
    17.50791, 17.27269, 17.1478, 17.23336, 17.82495, 17.98757, 17.42439,
    17.01356, 16.21792,
  12.11701, 12.14221, 12.17525, 12.19397, 12.17715, 12.16672, 12.17922,
    12.18891, 12.23183, 12.25685, 12.95835, 12.92408, 12.25749, 12.4347,
    12.5079, 12.26838, 12.211, 12.23046, 12.23461, 12.64642, 12.8016,
    12.43998, 12.42649, 12.84992, 13.0041, 12.62909, 14.83481, 16.00706,
    13.87928, 12.72252,
  12.44374, 12.40189, 12.29309, 12.48638, 12.32872, 12.2137, 12.25095,
    12.28616, 12.34011, 12.4603, 12.83549, 13.2731, 13.48992, 12.9257,
    12.77274, 12.72988, 12.34409, 12.35317, 12.69823, 13.06834, 13.01278,
    12.52161, 12.5244, 13.03284, 16.54814, 16.63275, 15.91326, 18.42941,
    14.76275, 13.23848,
  12.38363, 12.35878, 12.31988, 12.37705, 12.30142, 12.24398, 12.25897,
    12.31239, 12.40027, 12.44461, 12.50815, 12.89235, 13.16723, 13.54573,
    13.53434, 12.82543, 12.76932, 13.00177, 12.9711, 13.05112, 13.55946,
    14.53432, 15.39711, 14.86124, 19.37461, 21.33154, 17.91352, 18.13649,
    14.60101, 13.64684,
  12.31456, 12.29615, 12.44323, 12.54686, 12.73918, 13.09989, 13.10897,
    12.88962, 12.94653, 13.17604, 13.19734, 13.46714, 13.24771, 13.11168,
    13.88541, 14.59857, 13.92724, 13.07405, 13.06926, 13.1786, 15.29318,
    16.38725, 15.76767, 19.76717, 20.95584, 19.31331, 20.47603, 17.79462,
    14.55807, 13.09505,
  12.60088, 12.41978, 12.6058, 12.9021, 13.17244, 13.31496, 13.2841,
    13.13284, 13.67951, 14.02744, 13.84435, 13.58559, 13.32784, 13.51424,
    14.14912, 14.60378, 13.64716, 13.01269, 13.32183, 17.51151, 18.48414,
    14.96058, 14.92334, 16.99374, 18.46477, 18.1499, 17.51928, 18.02202,
    18.28803, 14.30569,
  12.59117, 12.62559, 13.30655, 14.24595, 14.14246, 13.63991, 13.69186,
    13.50949, 13.27837, 13.35017, 13.20742, 14.74448, 16.26157, 16.36086,
    15.57816, 21.61497, 26.59961, 19.89275, 15.83602, 18.09729, 16.6245,
    13.85737, 14.41266, 14.99151, 17.51998, 16.85261, 19.56385, 30.34188,
    26.29693, 13.81863,
  12.69846, 12.97353, 13.7682, 14.68752, 14.75667, 14.26057, 14.85205,
    16.30178, 16.54935, 16.45637, 17.11759, 16.84981, 16.02797, 15.93389,
    20.51026, 27.11624, 25.18692, 18.24204, 16.04407, 15.79429, 14.54636,
    13.84209, 14.32448, 16.30412, 17.64985, 15.41241, 24.59631, 37.70045,
    26.29476, 12.61092,
  12.88818, 13.20406, 14.13699, 14.97535, 14.84845, 16.59675, 18.39459,
    16.93132, 16.03525, 16.27611, 16.42287, 15.40841, 14.47311, 14.5827,
    17.26928, 19.10737, 17.68586, 15.99664, 14.81449, 14.53761, 14.05679,
    13.89848, 14.94489, 17.01354, 16.85302, 15.06331, 27.96525, 32.20967,
    18.05848, 12.78488,
  14.29721, 14.51108, 15.72404, 15.78181, 16.26114, 18.14389, 17.40177,
    15.85189, 15.93081, 16.22496, 15.7976, 14.85674, 14.33193, 17.44289,
    18.85999, 16.23122, 16.3611, 17.56596, 17.40895, 15.40007, 13.83452,
    14.96801, 18.50303, 19.00818, 16.37715, 16.4113, 23.3525, 22.04173,
    14.58974, 12.86892,
  16.60549, 17.85589, 19.62448, 20.70547, 20.88633, 18.18574, 15.30061,
    15.16282, 15.08834, 14.58397, 15.87666, 18.88882, 19.96242, 19.67847,
    18.77183, 18.65341, 19.25656, 19.78237, 18.89466, 17.61249, 17.38712,
    18.31136, 19.54073, 18.06524, 22.30403, 30.15907, 24.5861, 15.79552,
    13.46498, 12.34008,
  25.77778, 28.84795, 26.51492, 22.05167, 21.39351, 20.36012, 17.7967,
    19.42166, 20.74476, 27.01562, 29.48386, 20.50126, 17.86451, 17.21996,
    16.58797, 17.56578, 18.8796, 18.95632, 17.91129, 17.885, 20.11046,
    20.1661, 17.52261, 15.58057, 19.60947, 23.81734, 18.3689, 13.18817,
    12.60127, 12.19531,
  37.20757, 29.50283, 30.51902, 30.6997, 29.25052, 26.05397, 28.73706,
    26.6714, 22.21004, 26.78415, 26.19427, 16.12865, 16.83065, 17.69085,
    16.7081, 17.102, 16.92695, 16.94852, 16.49356, 17.12624, 19.93476,
    18.97872, 15.29868, 18.47912, 19.90006, 14.84032, 12.64991, 12.85298,
    12.76141, 12.32172,
  42.06897, 38.52677, 52.61045, 58.05249, 57.44957, 50.41957, 38.51646,
    25.54544, 23.34983, 22.19629, 19.00286, 14.42613, 18.94203, 21.01613,
    17.80047, 17.17596, 17.4787, 16.79965, 16.27604, 18.62247, 20.26109,
    17.54873, 14.895, 20.12381, 20.93921, 14.10365, 12.73202, 13.00174,
    13.2225, 12.55089,
  50.18657, 71.50313, 74.05263, 71.25262, 63.70177, 54.11904, 43.7531,
    38.84629, 30.82694, 27.62935, 32.5348, 32.65237, 36.27954, 36.38418,
    30.29668, 22.29801, 17.92334, 19.21288, 20.53855, 21.77002, 19.48148,
    18.91841, 20.32046, 17.58723, 15.21519, 13.32207, 12.80419, 12.65485,
    13.05406, 12.55935,
  38.17398, 46.70689, 46.06862, 44.31724, 38.62211, 40.40669, 53.7283,
    52.49828, 43.22563, 44.68506, 44.34011, 33.57957, 26.6803, 31.82896,
    32.48599, 21.48863, 20.80602, 20.96368, 22.92513, 24.32831, 22.31452,
    19.77217, 17.32126, 14.36918, 12.97528, 13.32084, 12.88949, 12.56538,
    12.59662, 12.3473,
  27.89984, 28.25957, 28.12254, 27.08213, 25.87897, 30.53189, 37.97917,
    35.83751, 33.15516, 33.49557, 30.28132, 22.82239, 18.79577, 22.87295,
    22.83907, 20.29182, 21.76371, 20.28932, 20.89716, 21.0663, 18.05963,
    15.70292, 13.50665, 13.35097, 13.49353, 13.24571, 12.91964, 12.62751,
    12.50171, 12.27624,
  26.01786, 25.24524, 23.97721, 23.12239, 23.61518, 24.69803, 25.35335,
    25.02453, 24.32749, 22.94406, 19.46079, 19.65894, 22.27481, 20.98693,
    20.30159, 20.38911, 20.16521, 18.4246, 19.4115, 18.32254, 13.99127,
    14.07196, 13.8524, 13.51154, 13.32087, 13.24614, 12.82774, 12.44465,
    12.43536, 12.27021,
  23.08296, 22.21237, 21.27706, 21.60402, 22.1524, 22.9649, 23.43875,
    23.45119, 22.55309, 19.91136, 19.33859, 22.40722, 23.36147, 22.88978,
    24.17586, 22.36687, 18.85275, 16.58328, 18.63818, 17.35419, 14.00624,
    14.22255, 14.0906, 13.66028, 12.95686, 12.99321, 12.71843, 12.30733,
    12.28856, 12.20777,
  22.56464, 22.32702, 21.10558, 20.88794, 21.31726, 21.59066, 21.71758,
    21.40596, 19.96641, 18.55939, 20.77435, 21.81147, 19.42303, 20.26974,
    20.98002, 19.7964, 19.03861, 18.88568, 20.52454, 19.45135, 16.5436,
    14.95186, 14.125, 13.6788, 12.8241, 12.69248, 12.59282, 12.31016,
    12.24374, 12.18879,
  23.01007, 22.98512, 21.55794, 20.49133, 20.65922, 20.56752, 20.35809,
    19.9069, 19.05334, 20.39418, 21.53187, 18.84266, 17.09434, 17.19811,
    16.89817, 16.3893, 17.47323, 19.11685, 20.18176, 20.45663, 19.17347,
    16.40734, 14.20717, 13.73394, 13.10998, 12.69636, 12.53892, 12.33081,
    12.25558, 12.19353,
  22.69886, 22.88441, 21.50733, 20.30363, 20.09251, 20.04501, 19.89995,
    19.5778, 19.61944, 21.32827, 19.87503, 16.34196, 16.53176, 16.48605,
    15.77406, 15.29912, 15.70521, 16.4526, 17.15608, 17.31532, 17.67531,
    17.26794, 15.56334, 14.26642, 13.4889, 12.90899, 12.53515, 12.32732,
    12.26389, 12.19451,
  23.25158, 22.6558, 21.2884, 20.43677, 20.17736, 19.81338, 19.88371,
    19.65476, 20.28881, 20.60679, 17.50257, 15.00604, 15.58245, 15.6772,
    15.34176, 15.18687, 14.93438, 14.79472, 15.10141, 15.08591, 16.234,
    16.29979, 15.62872, 15.91623, 14.73961, 13.20546, 12.63138, 12.40317,
    12.2731, 12.19914,
  23.39425, 22.8044, 21.03488, 20.25372, 20.7, 20.97587, 20.87535, 19.97074,
    20.13149, 18.94635, 15.68389, 14.52775, 14.93378, 15.13695, 14.89375,
    15.08698, 14.83879, 14.16042, 14.12341, 14.19064, 15.31382, 14.96123,
    14.02447, 15.58062, 15.80931, 13.86019, 12.85939, 12.79569, 12.50147,
    12.22433,
  23.01231, 22.58362, 21.61061, 21.37233, 21.64964, 21.89186, 22.20658,
    21.74515, 21.3547, 18.28652, 15.08205, 14.92545, 15.44964, 15.84962,
    15.5228, 15.39952, 15.42667, 14.74763, 14.14015, 14.24287, 14.42398,
    14.06538, 13.64827, 14.03327, 14.98452, 15.26003, 14.11309, 13.14286,
    12.83765, 12.32547,
  23.11382, 23.63486, 21.7925, 21.24893, 21.76687, 21.82651, 21.43846,
    21.19996, 21.68394, 18.55901, 15.17231, 15.24292, 15.71877, 15.99913,
    15.92588, 15.81793, 15.50004, 15.18816, 14.61195, 14.15999, 14.09736,
    14.005, 13.93628, 13.54366, 13.56011, 14.90868, 15.02564, 13.8193,
    13.6438, 12.65132,
  23.49105, 25.37965, 23.91151, 22.32774, 21.72929, 21.09241, 21.55978,
    22.21917, 21.04018, 17.94545, 15.69618, 15.71415, 16.11226, 15.87808,
    15.44839, 15.44531, 15.1549, 15.07251, 14.85737, 14.33879, 14.38218,
    14.3407, 13.69634, 13.29613, 13.33479, 13.99502, 15.33172, 14.44631,
    13.7019, 12.64003,
  24.44017, 26.38485, 23.99578, 22.00009, 21.13181, 20.36168, 21.95766,
    22.53329, 19.5948, 16.87376, 16.05767, 15.97332, 15.96494, 15.62732,
    15.27903, 15.09361, 14.84057, 14.95556, 14.82007, 14.31971, 14.47892,
    15.24834, 15.18902, 14.74156, 14.7856, 14.89969, 16.68758, 16.15219,
    13.56691, 12.23243,
  24.43454, 25.07011, 22.57365, 21.41998, 21.65366, 21.30124, 22.21843,
    21.08948, 17.79383, 16.28692, 15.7363, 15.56991, 15.46309, 15.49209,
    15.76084, 15.43032, 14.85353, 14.81291, 15.25603, 15.66507, 16.00167,
    15.88326, 15.45845, 15.11917, 15.36757, 15.33331, 15.96432, 17.7498,
    15.94154, 12.76769,
  22.30696, 21.29461, 21.41801, 22.5797, 23.28145, 23.79966, 22.9305,
    19.63538, 17.05595, 16.06997, 14.91471, 14.40992, 14.55945, 14.89054,
    15.4667, 15.66394, 15.70811, 16.09729, 15.93066, 15.64409, 15.69871,
    15.18997, 14.27976, 13.94341, 14.26716, 14.6735, 14.7692, 15.015,
    15.63843, 13.24509,
  21.222, 21.10641, 21.42835, 21.84384, 22.14102, 23.71108, 23.48211,
    19.4269, 16.63977, 16.00506, 15.52561, 15.82059, 16.40268, 16.40537,
    16.40264, 16.58699, 15.94946, 15.29148, 15.02758, 14.38855, 13.97517,
    13.84508, 13.53212, 13.37914, 13.46328, 14.00901, 14.168, 13.59696,
    13.24454, 12.43614,
  10.84216, 10.86247, 10.89296, 10.90699, 10.89918, 10.89234, 10.89627,
    10.90314, 10.93661, 10.93443, 11.59956, 11.57738, 10.95033, 11.11633,
    11.18668, 10.98177, 10.93734, 10.94541, 10.93054, 11.3596, 11.51256,
    11.14235, 11.11328, 11.50594, 11.57757, 11.16571, 13.14146, 14.26369,
    12.53223, 11.46933,
  11.1324, 11.0973, 11.0013, 11.18177, 11.04982, 10.93636, 10.95966,
    10.98842, 11.03425, 11.13074, 11.55751, 11.95413, 12.06853, 11.57328,
    11.44456, 11.39456, 11.04418, 11.057, 11.37801, 11.8072, 11.76718,
    11.20438, 11.15606, 11.62437, 14.83588, 14.85313, 14.53517, 17.18074,
    13.71107, 12.09126,
  11.11445, 11.09552, 11.05758, 11.11597, 11.02578, 10.93791, 10.94654,
    11.00731, 11.08306, 11.13313, 11.18765, 11.5593, 11.84832, 12.10804,
    12.09307, 11.48269, 11.40784, 11.63084, 11.6395, 11.68512, 12.0805,
    12.94466, 13.6832, 13.04599, 17.61767, 19.75261, 16.59637, 17.06886,
    13.57167, 12.51405,
  11.03235, 11.0083, 11.13849, 11.21092, 11.36518, 11.67593, 11.68217,
    11.48199, 11.50309, 11.71679, 11.77623, 12.0443, 11.82299, 11.69567,
    12.41609, 13.053, 12.43158, 11.63276, 11.56456, 11.55848, 13.60888,
    14.72307, 14.09187, 17.801, 19.22499, 18.20386, 19.47835, 16.69851,
    13.36762, 11.90132,
  11.28986, 11.09279, 11.25746, 11.49322, 11.74029, 11.90333, 11.86243,
    11.69591, 12.18334, 12.61571, 12.53058, 12.21173, 11.88116, 12.02623,
    12.66211, 13.06169, 11.96588, 11.30281, 11.56725, 15.45471, 16.58578,
    13.46847, 13.4042, 15.70343, 17.15887, 16.82053, 16.42771, 16.71412,
    16.73326, 12.92488,
  11.24731, 11.21169, 11.81849, 12.66487, 12.63533, 12.20667, 12.22007,
    12.04133, 11.86835, 12.00281, 11.81038, 13.06673, 14.38604, 14.48458,
    13.5968, 18.77233, 23.25903, 17.47642, 13.90497, 16.46298, 15.2271,
    12.47765, 13.09828, 13.6577, 16.19121, 15.53064, 17.48369, 27.76052,
    24.60325, 12.55754,
  11.2595, 11.50599, 12.26385, 13.14244, 13.32209, 12.7786, 13.12476,
    14.45315, 14.62584, 14.50023, 15.05763, 14.8985, 14.1885, 13.96163,
    18.06625, 24.54856, 23.23645, 16.59764, 14.47413, 14.43189, 13.2788,
    12.55504, 13.00386, 14.88141, 16.29663, 13.97992, 22.48103, 36.11668,
    25.55501, 11.33042,
  11.40767, 11.69529, 12.59804, 13.38585, 13.19934, 14.70896, 16.46571,
    15.24662, 14.35494, 14.51097, 14.63864, 13.60798, 12.61337, 12.60071,
    15.51035, 17.71266, 16.19919, 14.42658, 13.44396, 13.24908, 12.80969,
    12.61064, 13.54963, 15.60291, 15.51074, 13.58214, 26.50356, 31.56334,
    17.07495, 11.46204,
  12.52008, 12.66515, 13.80152, 13.85595, 14.19333, 16.3518, 15.88153,
    14.09644, 14.11742, 14.3615, 13.80974, 12.85099, 12.36082, 15.52509,
    17.10504, 14.67899, 14.8738, 16.05633, 15.89157, 14.0232, 12.49733,
    13.50483, 16.91561, 17.55941, 15.03816, 14.89616, 22.21113, 21.06077,
    13.10198, 11.59972,
  14.32018, 15.37131, 17.09051, 18.22886, 18.5484, 16.1475, 13.35779,
    13.12409, 13.17691, 12.65115, 13.75082, 16.60179, 17.91688, 18.06469,
    17.35924, 17.07671, 17.58991, 18.1942, 17.52318, 16.33569, 15.94274,
    16.82809, 18.21848, 16.92115, 20.56045, 28.04134, 23.16717, 14.61278,
    12.20212, 11.07256,
  21.49537, 24.3303, 22.83305, 19.02342, 18.63929, 17.68336, 15.27298,
    16.9963, 18.19048, 23.90803, 26.40384, 18.69773, 16.60538, 15.99157,
    15.23472, 16.29216, 17.58975, 17.649, 16.68464, 16.68521, 18.84418,
    18.88964, 16.31545, 14.33154, 18.40143, 23.05318, 17.66141, 11.98027,
    11.31369, 10.91151,
  31.20224, 24.76422, 25.68102, 25.5935, 24.2576, 21.65577, 24.68126,
    23.60455, 19.83302, 24.49924, 24.31917, 14.82532, 15.4021, 16.25206,
    15.41972, 15.81116, 15.63627, 15.66303, 15.19441, 15.79469, 18.69911,
    17.73722, 13.98642, 16.8656, 18.5722, 13.90366, 11.48272, 11.56494,
    11.48081, 11.04966,
  41.96664, 35.24341, 41.96729, 48.10627, 48.39857, 43.71891, 33.72121,
    22.24616, 20.8602, 20.23746, 17.27058, 12.9811, 17.38422, 19.48763,
    16.54509, 15.82404, 16.169, 15.48439, 14.86343, 17.25905, 19.02444,
    16.20047, 13.55956, 18.92322, 20.08347, 13.01211, 11.45542, 11.75388,
    11.9672, 11.30183,
  47.05423, 62.73176, 64.27415, 65.11072, 61.23177, 51.54025, 37.83696,
    34.06276, 27.21426, 24.63794, 29.52949, 30.07626, 33.92475, 33.99307,
    28.46324, 21.0654, 16.60175, 17.95141, 19.22388, 20.55957, 18.3298,
    17.5269, 19.09171, 16.79002, 14.32333, 12.0884, 11.54085, 11.40399,
    11.81711, 11.31845,
  32.64991, 40.33108, 41.29755, 41.89909, 37.26475, 37.16317, 47.75122,
    47.54292, 38.63207, 40.13034, 40.98651, 31.7941, 25.42897, 30.25198,
    31.02374, 20.25713, 19.51996, 19.66685, 21.42559, 22.96823, 20.97346,
    18.7207, 16.61341, 13.44073, 11.66173, 12.04206, 11.60937, 11.27645,
    11.32875, 11.09067,
  22.33235, 23.05773, 23.94973, 23.60815, 21.74226, 26.15429, 33.85804,
    31.43834, 29.49272, 31.01234, 28.74644, 21.49839, 17.3709, 21.57049,
    21.52072, 18.97698, 20.72367, 19.10911, 19.50327, 19.9544, 17.11089,
    14.82923, 12.50067, 12.21735, 12.23606, 11.94136, 11.63455, 11.35078,
    11.21468, 11.00176,
  21.18606, 20.75293, 19.90938, 19.01679, 19.09969, 20.22806, 21.00095,
    20.66879, 21.07063, 20.99723, 18.00405, 18.04115, 20.51158, 19.32467,
    18.89875, 19.2058, 19.22652, 17.41229, 18.1971, 17.32001, 12.94251,
    12.93971, 12.69347, 12.36581, 12.10178, 11.97127, 11.5638, 11.18471,
    11.14904, 10.9961,
  18.83861, 18.08044, 17.12406, 17.30598, 17.81906, 18.64498, 19.34318,
    19.9282, 19.71822, 17.71467, 17.06429, 20.29964, 21.75427, 21.37119,
    23.07341, 21.41485, 17.9708, 15.55797, 17.54723, 16.34832, 12.69572,
    12.90594, 12.8194, 12.43141, 11.73943, 11.72476, 11.46974, 11.04815,
    11.01686, 10.93793,
  18.46406, 18.12005, 16.7859, 16.56817, 17.07553, 17.53482, 17.98512,
    18.02908, 16.95144, 15.8839, 18.30463, 19.97074, 18.19343, 19.24228,
    20.25509, 19.06087, 18.04411, 17.5456, 19.08418, 17.90959, 14.95572,
    13.52248, 12.77066, 12.41279, 11.57075, 11.40936, 11.31813, 11.03637,
    10.97495, 10.92053,
  18.87659, 18.70787, 17.26101, 16.29257, 16.58113, 16.62201, 16.5701,
    16.28817, 15.71731, 17.44911, 19.33623, 17.49641, 16.02712, 16.27797,
    16.07622, 15.57903, 16.42787, 17.72819, 18.61818, 18.9111, 17.61739,
    14.96628, 12.83347, 12.44611, 11.85682, 11.41552, 11.25123, 11.05181,
    10.98205, 10.92227,
  18.46726, 18.63687, 17.36788, 16.25276, 16.14713, 16.06423, 15.85067,
    15.70142, 16.23972, 18.68128, 18.22613, 15.32267, 15.6201, 15.54983,
    14.78633, 14.23107, 14.44728, 15.04021, 15.70919, 16.01491, 16.47915,
    16.01639, 14.15814, 13.00883, 12.27024, 11.63452, 11.26328, 11.0542,
    10.99237, 10.92464,
  19.02896, 18.52041, 17.28777, 16.4318, 16.09818, 15.61626, 15.69876,
    15.906, 17.23093, 18.52578, 16.32095, 14.06192, 14.61709, 14.57575,
    14.15241, 13.93656, 13.68215, 13.57115, 13.91218, 13.86524, 15.04359,
    15.23488, 14.42967, 14.576, 13.34691, 11.90116, 11.34896, 11.12337,
    11.00351, 10.92648,
  19.29847, 18.74764, 17.04541, 16.12345, 16.44561, 16.70661, 16.89638,
    16.58698, 17.47685, 17.25278, 14.62321, 13.4678, 13.77511, 13.86145,
    13.61758, 13.89504, 13.73254, 13.04828, 12.92183, 12.93288, 14.1436,
    13.84984, 12.84303, 14.27682, 14.47823, 12.60274, 11.57582, 11.54768,
    11.24361, 10.94784,
  19.02411, 18.58084, 17.45914, 17.11586, 17.53762, 18.01364, 18.72116,
    18.83725, 18.9316, 16.43623, 13.77334, 13.65949, 14.09409, 14.48938,
    14.28631, 14.30272, 14.30243, 13.53036, 12.85266, 12.94267, 13.21427,
    12.86244, 12.38863, 12.80418, 13.79574, 14.0316, 12.86252, 11.92478,
    11.58938, 11.05458,
  18.9668, 19.10557, 17.59273, 17.32432, 18.08461, 18.49146, 18.44037,
    18.38713, 19.08451, 16.52452, 13.64397, 13.91143, 14.45877, 14.79447,
    14.79188, 14.70307, 14.30994, 13.91335, 13.30706, 12.88873, 12.81785,
    12.74664, 12.70646, 12.33801, 12.41814, 13.89188, 13.94619, 12.62336,
    12.41557, 11.41189,
  19.19009, 20.59492, 19.56478, 18.51909, 18.36589, 18.04729, 18.41372,
    18.94848, 18.0655, 15.8074, 14.06923, 14.39755, 14.93045, 14.73208,
    14.29061, 14.24615, 13.90571, 13.75996, 13.52034, 13.01353, 13.05087,
    13.06747, 12.45858, 12.06996, 12.14886, 12.89921, 14.24224, 13.29512,
    12.49126, 11.42771,
  20.21222, 21.85048, 20.24565, 18.72518, 17.89654, 17.05187, 18.60683,
    19.25996, 16.70857, 14.82488, 14.58109, 14.78983, 14.85441, 14.44572,
    13.99826, 13.79581, 13.56173, 13.59279, 13.43474, 12.96073, 13.1097,
    13.91952, 13.86382, 13.43856, 13.5589, 13.74821, 15.61402, 15.10084,
    12.39058, 10.99272,
  20.96515, 21.65694, 19.19956, 18.12924, 18.1652, 17.65044, 18.64656,
    17.86687, 15.17289, 14.43836, 14.46508, 14.4693, 14.27212, 14.13512,
    14.27818, 13.97924, 13.43582, 13.34307, 13.76347, 14.16521, 14.54253,
    14.5598, 14.23444, 13.92805, 14.23728, 14.32988, 15.05791, 16.88893,
    14.86161, 11.5113,
  19.47681, 18.36338, 18.17007, 19.26983, 19.71726, 19.8896, 19.18894,
    16.44812, 14.54458, 14.29548, 13.64286, 13.23271, 13.24228, 13.48451,
    14.00129, 14.15439, 14.15142, 14.44588, 14.37964, 14.23758, 14.36091,
    13.92896, 13.092, 12.78501, 13.15304, 13.66941, 13.82366, 14.15017,
    14.60864, 12.05157,
  18.36948, 17.98442, 18.35588, 18.87788, 19.07313, 20.27921, 19.8533,
    16.31738, 14.21051, 14.19417, 14.05268, 14.34505, 14.77186, 14.78982,
    14.88554, 15.04443, 14.44637, 13.84867, 13.60192, 13.034, 12.6721,
    12.60379, 12.31581, 12.17901, 12.30557, 12.9033, 13.13863, 12.49073,
    12.10482, 11.2299,
  9.467085, 9.48536, 9.519827, 9.533974, 9.526381, 9.516306, 9.522648,
    9.528828, 9.553441, 9.559355, 10.22486, 10.26182, 9.571901, 9.752356,
    9.854757, 9.635188, 9.578358, 9.57598, 9.551898, 9.977245, 10.184,
    9.82755, 9.79252, 10.15098, 10.20451, 9.779968, 11.79312, 13.20655,
    11.30855, 10.18193,
  9.750231, 9.750937, 9.62114, 9.829419, 9.701789, 9.565641, 9.587106,
    9.620323, 9.66256, 9.773684, 10.29111, 10.73695, 10.83431, 10.34705,
    10.14585, 10.11844, 9.703825, 9.67849, 10.01694, 10.54127, 10.52631,
    9.895766, 9.764008, 10.20178, 13.53523, 14.05254, 13.4068, 16.70582,
    12.71099, 10.92237,
  9.771594, 9.769139, 9.69004, 9.772958, 9.668083, 9.555859, 9.565988,
    9.643679, 9.730472, 9.801121, 9.869951, 10.31136, 10.71235, 10.95714,
    10.91976, 10.19691, 10.02566, 10.30389, 10.33874, 10.39278, 10.69011,
    11.45328, 12.20168, 11.48923, 16.60533, 20.00169, 15.82597, 16.78557,
    12.56957, 11.42134,
  9.666299, 9.647322, 9.777233, 9.829905, 9.962384, 10.32203, 10.37691,
    10.17358, 10.17729, 10.43568, 10.55396, 10.83426, 10.6033, 10.46667,
    11.24626, 11.85667, 11.25468, 10.36233, 10.19039, 10.01524, 11.9977,
    13.41387, 12.68287, 16.78137, 19.15055, 17.88223, 19.52495, 16.51258,
    12.49034, 10.76193,
  9.943911, 9.718523, 9.889833, 10.12655, 10.43023, 10.65025, 10.58744,
    10.37609, 10.87031, 11.51909, 11.54564, 11.11363, 10.62463, 10.75652,
    11.53055, 11.98828, 10.69549, 9.756349, 9.93927, 14.03734, 15.82407,
    12.22032, 12.03084, 14.88271, 16.64177, 16.14163, 16.23286, 16.29885,
    15.9812, 11.79778,
  9.886089, 9.784056, 10.41513, 11.41179, 11.51541, 11.00391, 10.93989,
    10.75886, 10.61398, 10.81077, 10.60268, 11.73105, 13.09302, 13.26389,
    12.41865, 17.14349, 22.08882, 16.35407, 12.39192, 15.48239, 14.59269,
    11.15287, 11.85676, 12.52912, 15.2356, 14.92822, 16.14894, 27.00027,
    24.84799, 11.62381,
  9.80928, 10.0558, 10.93273, 11.99208, 12.31482, 11.70963, 11.8653,
    13.12237, 13.2529, 13.1221, 13.63745, 13.66883, 13.02314, 12.66783,
    16.56078, 23.78441, 23.10675, 15.72649, 13.33348, 13.42957, 12.13172,
    11.31512, 11.80801, 13.86725, 15.57243, 12.96215, 21.62033, 38.0941,
    27.52129, 10.15904,
  9.936085, 10.25326, 11.2625, 12.19379, 12.0512, 13.49991, 15.32038,
    14.07157, 13.07231, 13.29817, 13.51507, 12.44707, 11.17888, 11.03933,
    14.1776, 17.05229, 15.37415, 13.32039, 12.29107, 12.09798, 11.63728,
    11.38518, 12.3368, 14.6354, 14.7063, 12.31678, 26.94538, 34.86492,
    17.36164, 10.22008,
  11.05882, 11.17432, 12.39219, 12.56418, 12.74592, 15.263, 14.98672,
    12.79407, 12.75815, 13.12059, 12.5468, 11.38143, 10.65326, 13.83749,
    15.89356, 13.41614, 13.62903, 15.08029, 14.84764, 12.92242, 11.22285,
    12.21918, 15.82504, 16.85739, 14.03953, 13.72205, 22.26745, 21.93115,
    11.94349, 10.41264,
  13.14711, 14.02092, 15.77773, 17.16694, 17.48132, 15.23106, 12.09454,
    11.72423, 11.81079, 11.12554, 12.03406, 15.19842, 16.67832, 17.00226,
    16.31378, 15.87834, 16.51453, 17.29984, 16.7129, 15.26444, 14.78174,
    15.89922, 17.63089, 16.29209, 19.5817, 27.78474, 23.23801, 13.86516,
    11.14669, 9.760143,
  19.01364, 22.55982, 22.0758, 18.239, 17.68143, 16.84726, 14.20884,
    15.90695, 16.80792, 22.60596, 26.14729, 17.91577, 15.71937, 15.04767,
    14.12614, 15.26927, 16.81746, 16.91993, 15.81474, 15.62179, 18.0731,
    18.40011, 15.68964, 13.31851, 17.83048, 23.46011, 17.80952, 10.90747,
    10.03957, 9.529259,
  33.97837, 26.97047, 24.19258, 24.27906, 22.86183, 19.97574, 23.56562,
    23.05903, 18.85327, 24.05606, 24.69461, 13.75016, 14.34594, 15.45012,
    14.47192, 15.09208, 14.84605, 14.79491, 14.29548, 14.90191, 18.18415,
    17.30791, 13.01405, 15.86732, 18.37266, 13.46093, 10.37204, 10.28404,
    10.19285, 9.707587,
  46.65451, 35.41777, 39.21328, 46.55322, 47.25008, 43.53527, 34.34328,
    21.46404, 20.15368, 19.98572, 17.11023, 11.55418, 16.54011, 19.18,
    15.77468, 15.12121, 15.41926, 14.65139, 14.00228, 16.70461, 18.82442,
    15.49428, 12.54407, 18.43442, 20.43945, 12.18883, 10.17592, 10.50569,
    10.75249, 10.02483,
  47.60692, 61.18661, 62.81955, 65.04876, 61.31219, 52.41998, 38.66318,
    34.32659, 27.37572, 23.12365, 28.45803, 29.18336, 33.2585, 33.53323,
    28.47137, 20.99117, 15.97954, 17.38036, 18.82696, 20.56917, 18.05626,
    16.97199, 19.28189, 16.71008, 13.82688, 10.9067, 10.27792, 10.14609,
    10.59937, 10.06436,
  31.0484, 38.47561, 40.42998, 42.3541, 38.32019, 37.42039, 47.77586,
    47.86346, 37.27263, 37.90753, 40.11013, 31.70418, 24.90019, 29.7776,
    31.6814, 20.10013, 19.1686, 19.29583, 21.19299, 23.48016, 21.66089,
    19.13808, 16.82209, 12.90825, 10.3741, 10.7824, 10.3319, 9.992106,
    10.0439, 9.781657,
  20.65033, 21.4664, 23.23853, 23.52439, 21.5411, 25.4635, 33.41388,
    30.59154, 28.08271, 30.06491, 28.66229, 21.54113, 16.89488, 21.55199,
    21.58235, 18.5658, 20.59308, 18.86045, 19.14695, 20.2494, 17.4692,
    14.72366, 11.71604, 11.21074, 11.0976, 10.71272, 10.37843, 10.11846,
    9.926692, 9.662655,
  19.98916, 19.8611, 19.26372, 18.2093, 17.88945, 19.09183, 20.21538,
    19.87596, 20.46067, 20.97137, 17.89079, 17.64264, 20.28185, 18.92692,
    18.5239, 18.95312, 19.2789, 17.24409, 17.84274, 17.36629, 12.24151,
    11.95279, 11.60747, 11.3593, 11.05223, 10.76242, 10.31357, 9.921489,
    9.845974, 9.656682,
  17.79339, 17.22491, 16.12749, 16.11664, 16.57386, 17.51229, 18.37656,
    19.04988, 18.94965, 17.12106, 16.31733, 19.87247, 21.70603, 20.94033,
    23.204, 21.57411, 17.97655, 15.09763, 17.19805, 16.25715, 11.75311,
    11.85239, 11.7067, 11.45517, 10.65872, 10.514, 10.23123, 9.713387,
    9.66434, 9.580847,
  17.52035, 17.19598, 15.61299, 15.23795, 15.74521, 16.32646, 16.84571,
    16.96065, 16.08598, 14.99983, 17.53453, 19.63162, 17.72102, 18.90069,
    20.55582, 19.29799, 17.97934, 16.93242, 18.57785, 17.31544, 13.85344,
    12.48976, 11.68623, 11.36531, 10.39053, 10.15395, 10.05568, 9.700094,
    9.614864, 9.549301,
  17.88586, 17.60598, 15.97751, 14.87337, 15.191, 15.27944, 15.32788,
    15.17501, 14.70586, 16.63377, 18.97408, 17.08862, 15.37334, 15.87838,
    15.94725, 15.41711, 16.17705, 17.26824, 17.96064, 18.29486, 16.92974,
    14.23829, 11.78754, 11.343, 10.65057, 10.11923, 9.942304, 9.711624,
    9.623242, 9.556425,
  17.25698, 17.33597, 15.96678, 14.80427, 14.73843, 14.74262, 14.61146,
    14.51976, 15.25722, 18.20641, 18.16115, 14.88988, 15.14085, 15.14215,
    14.34695, 13.5987, 13.69761, 14.19522, 14.89112, 15.56741, 16.23549,
    15.59504, 13.15371, 11.86236, 11.07029, 10.38632, 9.961967, 9.708876,
    9.616882, 9.555486,
  17.71628, 17.09704, 15.84882, 15.05024, 14.78004, 14.32365, 14.45509,
    14.80729, 16.57974, 18.48867, 16.34842, 13.69317, 14.21023, 14.08189,
    13.45775, 12.94009, 12.59026, 12.56138, 13.11777, 13.19368, 14.49713,
    14.76307, 13.47162, 13.62112, 12.35995, 10.73625, 10.04071, 9.80305,
    9.640373, 9.557379,
  17.98132, 17.3438, 15.72667, 14.83619, 15.22486, 15.54772, 15.85544,
    15.79768, 17.25438, 17.53782, 14.64962, 13.15985, 13.27496, 13.16495,
    12.65566, 12.80599, 12.77429, 12.19814, 12.09614, 12.02414, 13.37038,
    13.15915, 11.7771, 13.40819, 13.63224, 11.50326, 10.26205, 10.25647,
    9.922678, 9.587122,
  17.85237, 17.37818, 16.22523, 15.86683, 16.39668, 17.01578, 18.1422,
    18.79877, 19.23878, 16.72526, 13.64535, 13.26207, 13.42117, 13.66536,
    13.33157, 13.35155, 13.50995, 12.73326, 11.89196, 11.94208, 12.35208,
    11.9043, 11.21468, 11.73251, 12.86228, 12.9762, 11.65105, 10.7001,
    10.32324, 9.713716,
  17.77164, 17.67592, 16.30235, 16.20168, 17.30336, 18.08888, 18.3601,
    18.66771, 19.56749, 16.79005, 13.31702, 13.37139, 13.74397, 14.01715,
    13.94411, 13.87238, 13.519, 13.08759, 12.35752, 11.87989, 11.77203,
    11.62799, 11.62305, 11.22122, 11.2721, 12.80238, 12.9091, 11.53488,
    11.29792, 10.18859,
  17.93878, 18.93988, 18.40892, 17.88079, 17.98674, 18.05275, 18.64266,
    19.29622, 18.37892, 15.83925, 13.60011, 13.78443, 14.2368, 13.97761,
    13.42027, 13.37015, 13.00172, 12.83558, 12.5866, 11.96, 11.92271,
    11.93703, 11.35867, 10.88301, 10.86637, 11.67055, 13.18958, 12.30845,
    11.44499, 10.27525,
  18.99525, 20.30062, 19.52237, 18.53263, 17.73416, 17.03241, 18.88355,
    19.70432, 16.82771, 14.466, 14.06916, 14.24721, 14.24159, 13.66158,
    13.0734, 12.8371, 12.61275, 12.65865, 12.4862, 11.84955, 11.9508,
    12.83994, 12.86634, 12.33956, 12.3007, 12.51995, 14.63056, 14.24874,
    11.3248, 9.736085,
  20.29335, 20.86366, 18.56206, 17.96857, 18.02889, 17.56789, 18.68953,
    17.94962, 14.7968, 13.90399, 13.97375, 13.95057, 13.62259, 13.23383,
    13.30948, 13.02909, 12.44979, 12.3228, 12.71684, 13.08288, 13.47591,
    13.64649, 13.40328, 12.98132, 13.10355, 13.24914, 14.11819, 16.08347,
    14.06614, 10.31951,
  19.2815, 18.15672, 17.8875, 19.29386, 19.70574, 19.71118, 19.09649,
    16.14259, 13.96202, 13.89985, 13.23173, 12.61198, 12.35945, 12.46836,
    13.03676, 13.23973, 13.16062, 13.41499, 13.39132, 13.28027, 13.42204,
    12.97043, 12.07312, 11.66835, 12.01293, 12.60399, 12.81763, 13.30619,
    13.88847, 11.01687,
  18.3352, 17.92741, 18.21395, 18.71721, 18.86909, 20.10701, 19.71217,
    15.94588, 13.6916, 13.8705, 13.64465, 13.66981, 13.86285, 13.87291,
    13.98741, 14.12358, 13.52412, 12.89727, 12.60087, 11.98001, 11.57109,
    11.46698, 11.12121, 10.94509, 11.12047, 11.80556, 12.11722, 11.4584,
    11.02293, 9.990366,
  11.82008, 11.83432, 11.86781, 11.88601, 11.87621, 11.8696, 11.86803,
    11.87892, 11.90843, 11.91614, 12.59776, 12.72378, 11.91552, 12.06711,
    12.20989, 11.97845, 11.91236, 11.91929, 11.88526, 12.26424, 12.5397,
    12.22101, 12.20191, 12.53853, 12.5713, 12.12263, 14.00306, 15.73827,
    13.76416, 12.64309,
  12.04864, 12.08902, 11.93795, 12.16471, 12.06586, 11.91796, 11.93023,
    11.95614, 12.00353, 12.12027, 12.69602, 13.17792, 13.17663, 12.70884,
    12.45156, 12.48041, 12.04207, 11.98713, 12.30348, 12.87978, 12.94394,
    12.31088, 12.11217, 12.5775, 15.59291, 16.51508, 15.84141, 19.87132,
    15.3389, 13.50992,
  12.1004, 12.12353, 12.0336, 12.13749, 12.03106, 11.8985, 11.90526,
    11.98462, 12.07953, 12.1691, 12.25687, 12.69305, 13.1344, 13.35998,
    13.31634, 12.55355, 12.29567, 12.62404, 12.70447, 12.82087, 13.07084,
    13.78761, 14.48317, 13.81674, 18.37304, 22.53772, 18.41224, 19.88611,
    15.06502, 14.02622,
  12.02259, 12.00782, 12.14588, 12.1961, 12.29427, 12.68017, 12.75162,
    12.5281, 12.51763, 12.77473, 12.91181, 13.20301, 13.04367, 12.83401,
    13.6417, 14.23189, 13.73785, 12.76593, 12.54495, 12.2802, 14.20094,
    15.9173, 14.99478, 18.86555, 21.75925, 20.4025, 22.58801, 19.45716,
    14.96853, 13.26843,
  12.36008, 12.06816, 12.23463, 12.43128, 12.76364, 13.08524, 13.0161,
    12.73713, 13.18337, 13.95298, 14.06702, 13.59191, 12.97798, 13.03055,
    13.91442, 14.50435, 13.24096, 12.03481, 12.10875, 16.03938, 18.60611,
    14.64344, 14.24539, 17.18169, 19.37472, 18.90771, 19.15847, 19.12261,
    18.85423, 14.47392,
  12.28022, 12.09336, 12.69451, 13.72539, 13.91782, 13.39272, 13.26595,
    13.09234, 12.98462, 13.23168, 13.02836, 13.98525, 15.47557, 15.63366,
    14.90923, 18.66024, 24.09841, 19.12279, 14.60586, 17.79906, 17.32098,
    13.30809, 14.03172, 14.89853, 17.70209, 17.91046, 18.15439, 29.69515,
    29.20067, 14.42007,
  12.12455, 12.33224, 13.23827, 14.454, 14.78883, 14.07746, 14.08024,
    15.44164, 15.63756, 15.45496, 15.95777, 16.11902, 15.55014, 15.06606,
    18.5498, 25.90821, 25.88967, 18.39516, 15.64572, 15.86284, 14.43033,
    13.5046, 14.09918, 16.25495, 18.24449, 15.66176, 23.13197, 42.01684,
    33.42483, 12.75884,
  12.22879, 12.57537, 13.64433, 14.69625, 14.46446, 15.75614, 17.80993,
    16.66925, 15.50193, 15.72939, 16.03485, 15.0562, 13.51218, 13.21781,
    16.26772, 19.74623, 17.95859, 15.65334, 14.57666, 14.41812, 13.96501,
    13.69787, 14.76582, 17.26874, 17.4283, 14.72474, 29.56162, 41.25027,
    21.54321, 12.79194,
  13.3637, 13.52706, 14.72046, 14.97117, 15.055, 17.94568, 17.96797,
    15.31852, 15.16919, 15.65059, 15.08175, 13.71181, 12.75792, 15.87118,
    18.52636, 15.88977, 15.80841, 17.49007, 17.34524, 15.48698, 13.58008,
    14.602, 18.39677, 19.88755, 16.57172, 16.16088, 25.76945, 27.22965,
    14.59952, 13.00194,
  15.38552, 16.11888, 18.1144, 20.07434, 20.36941, 18.2975, 14.74251,
    14.21014, 14.24409, 13.62994, 14.19906, 17.31085, 18.92168, 19.59369,
    19.0139, 18.39125, 19.0315, 19.99103, 19.5917, 17.99559, 17.31931,
    18.43593, 20.47442, 19.17842, 21.91395, 31.29051, 27.77066, 17.07309,
    13.79769, 12.2063,
  20.68483, 25.19249, 25.13416, 20.78282, 20.41887, 19.97833, 17.0982,
    18.52356, 19.49613, 23.88201, 28.14563, 20.46357, 18.12116, 17.61067,
    16.63197, 17.82342, 19.65733, 19.88352, 18.77174, 18.27046, 20.83942,
    21.28055, 18.60235, 15.81626, 20.46554, 27.30961, 21.88085, 13.56057,
    12.51822, 11.90342,
  35.50952, 28.64249, 26.2538, 25.01013, 24.54062, 21.24038, 25.62072,
    26.10499, 21.27335, 25.9604, 27.28338, 16.03215, 16.48795, 17.93414,
    17.04975, 17.84564, 17.61848, 17.5897, 16.98556, 17.46742, 20.98828,
    20.35571, 15.62917, 18.19473, 21.67455, 16.84278, 13.03814, 12.69962,
    12.60193, 12.09186,
  47.83837, 33.83937, 37.35227, 44.77291, 48.35171, 46.72075, 39.10989,
    23.65744, 23.36235, 22.83965, 19.35479, 13.55094, 18.61864, 21.45848,
    18.48709, 17.93372, 18.20204, 17.28361, 16.48341, 19.32606, 21.87797,
    18.22956, 15.00404, 21.17334, 24.64546, 15.21579, 12.57721, 12.8976,
    13.11784, 12.45709,
  48.53734, 53.13674, 54.33167, 60.1906, 61.44633, 57.0963, 42.78908,
    36.77988, 30.61054, 24.36535, 29.43021, 30.44406, 35.03529, 35.64631,
    31.35752, 23.90509, 18.73545, 20.10221, 21.70162, 23.71823, 21.17025,
    19.26335, 22.4894, 20.57644, 17.3752, 13.44837, 12.65418, 12.56371,
    12.99321, 12.52966,
  32.12364, 36.26224, 40.96365, 48.97938, 51.14721, 45.88917, 48.07789,
    49.43249, 37.84341, 37.85019, 41.4273, 34.10543, 27.81995, 32.48784,
    34.74226, 23.2226, 22.14548, 22.30496, 24.23415, 26.54956, 24.473,
    22.30709, 20.60822, 16.48128, 12.86199, 13.21592, 12.74813, 12.41542,
    12.46026, 12.22125,
  21.80095, 24.58294, 29.74283, 32.85722, 30.85852, 29.38332, 33.805,
    31.09625, 28.19318, 31.24689, 30.90874, 23.9538, 19.21391, 24.56674,
    24.74837, 21.52564, 23.88524, 22.07371, 21.96509, 23.49218, 20.69504,
    18.20828, 14.91825, 13.93627, 13.61531, 13.20798, 12.8065, 12.54582,
    12.33504, 12.07348,
  20.18779, 21.31371, 21.69291, 20.20347, 18.41571, 19.07697, 20.63179,
    19.91585, 20.72981, 22.10485, 19.16735, 18.90878, 22.30929, 21.40244,
    21.3513, 21.826, 22.56963, 20.47756, 20.74837, 21.14202, 15.46335,
    14.92128, 14.27519, 13.9307, 13.62832, 13.25927, 12.74216, 12.35523,
    12.24055, 12.05826,
  17.29546, 17.05287, 15.66907, 14.99897, 15.24392, 16.60714, 17.65877,
    18.31802, 18.60157, 17.01719, 16.42773, 20.80943, 23.53905, 22.83958,
    26.16293, 24.92927, 21.31299, 18.12407, 20.35805, 20.03923, 14.63198,
    14.60053, 14.25905, 14.05785, 13.21301, 12.9772, 12.70994, 12.13689,
    12.06404, 11.98066,
  16.62905, 16.1491, 14.32397, 13.80833, 14.35679, 15.03805, 15.72699,
    16.02595, 15.2865, 14.14711, 17.24606, 20.58215, 19.02128, 20.83391,
    23.57855, 22.59837, 21.40464, 20.11585, 21.99671, 20.81161, 16.59729,
    15.13223, 14.27877, 14.00002, 12.9076, 12.59775, 12.52778, 12.12164,
    12.02021, 11.94656,
  16.72952, 16.1185, 14.43866, 13.25647, 13.64018, 13.86107, 14.1023,
    14.0503, 13.42488, 15.50399, 18.90696, 17.74523, 16.46956, 17.95791,
    18.7397, 18.49485, 19.58515, 20.85876, 21.29856, 21.54706, 19.92999,
    17.18468, 14.41477, 13.93155, 13.16746, 12.55034, 12.38419, 12.14701,
    12.0231, 11.95094,
  15.90862, 15.72742, 14.39654, 13.25082, 13.28645, 13.45611, 13.36666,
    13.11804, 13.77804, 17.21353, 18.23582, 15.32787, 16.43984, 17.37796,
    17.14696, 16.66462, 16.93801, 17.42929, 17.81523, 18.61105, 19.42719,
    18.7699, 15.83333, 14.45202, 13.57789, 12.87566, 12.40308, 12.13451,
    12.0195, 11.95258,
  16.47764, 15.55714, 14.40627, 13.67799, 13.5438, 13.04888, 13.03198,
    13.24135, 15.2414, 17.81171, 16.29635, 14.18334, 15.79607, 16.48946,
    16.33716, 15.97778, 15.57978, 15.36008, 15.90262, 16.08828, 17.46051,
    18.0531, 16.14684, 16.32893, 15.01109, 13.29629, 12.47695, 12.23126,
    12.03967, 11.94771,
  16.9022, 15.99641, 14.47793, 13.55601, 13.94144, 14.10201, 14.33645,
    14.28393, 16.11339, 17.12352, 14.55818, 13.84779, 14.98899, 15.6068,
    15.45062, 15.68651, 15.64799, 15.00732, 14.88989, 14.75384, 16.20191,
    16.37744, 14.39664, 16.13985, 16.37107, 14.09784, 12.63601, 12.68532,
    12.34626, 11.98777,
  16.89356, 16.14206, 15.05117, 14.55569, 14.98445, 15.46945, 16.81718,
    17.7893, 18.53827, 16.43428, 13.54535, 14.07339, 15.1435, 16.06366,
    16.02523, 16.13458, 16.41459, 15.63303, 14.61719, 14.60603, 15.20522,
    14.77694, 13.76859, 14.34541, 15.47863, 15.58443, 14.18984, 13.15548,
    12.77657, 12.14288,
  16.77182, 16.50059, 15.04088, 14.7583, 15.82181, 16.81762, 17.4593,
    18.04265, 19.17479, 16.734, 13.32413, 14.22571, 15.38471, 16.35483,
    16.66736, 16.84115, 16.55729, 16.01294, 15.08833, 14.55373, 14.50453,
    14.25189, 14.21907, 13.81303, 13.79334, 15.40704, 15.57066, 14.04838,
    13.75511, 12.71253,
  16.94733, 17.70735, 17.00268, 16.3551, 16.66697, 17.1194, 18.01913,
    18.8849, 18.06431, 15.78744, 13.57109, 14.50545, 15.85028, 16.37961,
    16.26066, 16.42621, 15.98485, 15.6247, 15.34585, 14.59659, 14.54136,
    14.61465, 13.98731, 13.36735, 13.29275, 14.19477, 15.69347, 14.91234,
    13.89606, 12.81521,
  18.03276, 19.00228, 18.1799, 17.16967, 16.70685, 16.26605, 18.52649,
    19.66812, 16.5157, 14.08325, 13.96548, 15.00798, 16.0464, 16.184,
    15.91232, 15.71765, 15.3716, 15.31436, 15.154, 14.41994, 14.51453,
    15.47453, 15.46583, 14.7843, 14.75011, 15.00522, 17.14133, 16.99265,
    13.83581, 12.1725,
  19.4349, 20.00813, 17.3696, 16.88524, 17.23543, 17.01597, 18.50965,
    17.96717, 14.29397, 13.31946, 13.93764, 14.89816, 15.53759, 15.75479,
    16.11927, 15.85647, 15.13702, 14.86421, 15.16741, 15.49111, 15.99744,
    16.42898, 16.12851, 15.58374, 15.68883, 15.87894, 16.78514, 18.78977,
    16.86109, 12.85684,
  18.40132, 17.18413, 16.91184, 18.86164, 19.43048, 19.45325, 19.00371,
    15.824, 13.17323, 13.32383, 13.28269, 13.54048, 14.15547, 14.87945,
    15.8326, 16.05954, 15.80532, 15.95713, 15.87321, 15.76758, 16.07616,
    15.74767, 14.7601, 14.24791, 14.63529, 15.26172, 15.51421, 16.05274,
    16.64459, 13.73279,
  17.68913, 17.23341, 17.85773, 18.82208, 19.0546, 20.13462, 19.61183,
    15.47873, 12.95663, 13.46935, 13.75508, 14.51934, 15.52847, 16.2459,
    16.74211, 16.90966, 16.24414, 15.53964, 15.16257, 14.53145, 14.14268,
    14.01948, 13.68577, 13.48922, 13.70247, 14.40913, 14.73188, 14.02581,
    13.581, 12.51943,
  12.20887, 12.24106, 12.26808, 12.28617, 12.27701, 12.26709, 12.27147,
    12.28051, 12.30048, 12.33673, 13.13317, 13.38213, 12.34885, 12.53883,
    12.75258, 12.41655, 12.31033, 12.33401, 12.32475, 12.80442, 13.23339,
    12.84447, 12.81608, 13.21411, 13.26348, 12.74885, 14.90117, 17.43694,
    14.8194, 13.35402,
  12.48665, 12.57632, 12.3618, 12.64684, 12.50274, 12.30345, 12.33665,
    12.36809, 12.4274, 12.61292, 13.25689, 13.86646, 13.96062, 13.4361,
    13.0197, 13.06956, 12.47027, 12.42283, 12.88884, 13.65728, 13.71465,
    12.91276, 12.64743, 13.33547, 17.02017, 19.08177, 17.61717, 23.17484,
    16.86842, 14.47829,
  12.53958, 12.58034, 12.48248, 12.59411, 12.44843, 12.29425, 12.30209,
    12.40236, 12.52695, 12.64435, 12.78145, 13.3014, 13.82692, 14.17156,
    14.17639, 13.13346, 12.83849, 13.33151, 13.42514, 13.58536, 13.9081,
    14.89487, 15.84674, 15.3003, 20.63313, 26.94298, 21.3132, 23.42077,
    16.55188, 15.27295,
  12.48162, 12.46416, 12.63579, 12.7331, 12.8238, 13.26607, 13.3757,
    13.11219, 13.07569, 13.37068, 13.62161, 13.96826, 13.80494, 13.47405,
    14.51973, 15.37182, 14.87221, 13.55017, 13.17688, 12.91861, 15.37228,
    17.80054, 16.59359, 21.39187, 25.44976, 23.28002, 27.08981, 22.53024,
    16.41045, 14.27269,
  12.9377, 12.53566, 12.76629, 13.00599, 13.40827, 13.75041, 13.61844,
    13.32027, 13.86998, 15.05501, 15.42486, 14.55236, 13.56744, 13.86775,
    15.06821, 15.59226, 14.09513, 12.48864, 12.71212, 17.48411, 21.24068,
    16.08803, 15.60919, 18.98318, 21.60233, 21.06551, 21.71653, 22.24293,
    21.93293, 15.76695,
  12.79445, 12.58544, 13.34159, 14.60927, 14.99377, 14.34834, 13.89278,
    13.71607, 13.61235, 14.04656, 13.95057, 14.9727, 17.01997, 17.31775,
    16.77868, 21.2596, 28.41565, 22.04164, 16.08063, 19.80352, 19.3736,
    14.27611, 15.13875, 16.3476, 19.28279, 19.74211, 19.54195, 33.33809,
    34.50523, 15.72708,
  12.61138, 12.90333, 14.01513, 15.50605, 16.09749, 15.30353, 14.94772,
    16.79452, 17.29948, 17.17205, 17.85313, 18.08839, 17.23214, 16.76638,
    21.10791, 30.20858, 29.81654, 20.41504, 17.18904, 17.51736, 15.67264,
    14.38167, 15.13981, 17.78666, 20.11239, 17.39314, 24.06209, 45.00059,
    38.84227, 13.77376,
  12.70604, 13.1764, 14.50491, 15.86718, 15.65492, 17.14031, 19.84152,
    18.5473, 16.95565, 17.38358, 17.70944, 16.60484, 14.61096, 14.44485,
    18.2153, 22.4115, 19.71267, 17.12841, 15.76267, 15.5164, 14.88291,
    14.52958, 15.90989, 19.03773, 19.25322, 16.40046, 31.25823, 45.9304,
    24.01958, 13.64879,
  14.16602, 14.43022, 15.68752, 16.0328, 16.37889, 20.29692, 20.51231,
    16.76981, 16.67661, 17.26992, 16.56643, 14.7709, 13.628, 17.338,
    21.13203, 17.84104, 17.07647, 19.11115, 19.04189, 16.89006, 14.44271,
    15.73974, 20.27998, 22.42961, 18.18373, 17.88358, 28.25822, 31.19361,
    16.0613, 13.74674,
  16.50146, 17.05175, 19.61718, 22.97546, 23.03387, 20.5968, 16.04572,
    15.24044, 15.276, 14.63487, 15.123, 19.04922, 21.04993, 21.78496,
    20.91859, 20.09964, 21.00329, 22.1222, 21.46244, 19.47656, 18.88823,
    20.20404, 22.55277, 21.34498, 24.52872, 36.3362, 33.20652, 19.02905,
    14.63241, 12.71114,
  23.52068, 30.64741, 31.08097, 23.29469, 22.99362, 22.5861, 19.83665,
    21.13364, 22.36411, 26.12439, 32.17741, 23.57616, 20.30067, 19.55993,
    18.38855, 19.78459, 22.2191, 22.53967, 21.06293, 19.75599, 22.76151,
    23.35869, 20.25792, 17.07385, 22.37443, 30.62446, 24.85749, 14.31308,
    13.14087, 12.29239,
  41.53899, 34.56565, 30.40934, 26.68283, 27.36663, 22.67611, 27.40554,
    28.17502, 23.71958, 28.85725, 30.52159, 17.46357, 18.3848, 20.11509,
    18.94874, 20.08326, 19.94671, 19.94437, 19.03421, 19.22576, 23.22303,
    22.35236, 16.65026, 19.65806, 24.74876, 19.02397, 13.97854, 13.33447,
    13.21225, 12.54701,
  55.54279, 41.66972, 43.76203, 50.53552, 52.79464, 49.93245, 44.35527,
    37.90645, 44.18103, 31.16758, 21.06758, 15.87107, 22.08414, 24.21837,
    21.51075, 20.0041, 20.61154, 19.52211, 18.17277, 21.51397, 24.7592,
    19.7739, 15.95909, 23.1616, 28.63888, 16.59858, 13.18644, 13.55978,
    13.81479, 13.0437,
  62.37083, 52.80597, 56.4241, 62.7375, 65.89132, 66.30505, 58.98834,
    58.21395, 48.05751, 30.96942, 34.721, 37.45204, 42.7904, 43.52002,
    38.14014, 27.38035, 21.18405, 23.0023, 25.20198, 27.76149, 24.54205,
    20.83464, 25.29904, 23.18632, 19.36855, 14.28578, 13.26196, 13.12684,
    13.61226, 13.14298,
  47.40604, 59.31194, 68.61896, 75.63209, 76.45933, 67.47026, 66.19381,
    68.29429, 46.36478, 45.60231, 52.11835, 43.10053, 34.86663, 41.52793,
    42.76838, 28.01364, 25.97097, 26.44368, 28.72297, 30.95912, 27.0389,
    24.92024, 23.38417, 18.30217, 13.46459, 13.81312, 13.33161, 12.9673,
    12.9882, 12.73376,
  34.85776, 45.86493, 52.80127, 52.27154, 46.07896, 45.32644, 48.99612,
    39.51424, 38.34939, 44.3571, 40.58337, 31.27583, 25.19104, 31.2897,
    30.16199, 25.79068, 28.55332, 26.20885, 24.86908, 26.4087, 22.53679,
    20.10708, 16.64392, 15.05664, 14.33276, 13.83282, 13.35296, 13.10156,
    12.85347, 12.53753,
  27.74525, 29.57965, 29.9948, 26.584, 24.00937, 27.40716, 29.52086,
    26.17019, 30.05906, 32.0708, 25.15424, 24.04255, 27.95838, 25.63758,
    25.47098, 25.76458, 26.96534, 23.79056, 22.97484, 24.46518, 17.08348,
    16.17892, 15.35242, 15.02421, 14.58231, 13.95354, 13.31426, 12.8654,
    12.71014, 12.50504,
  22.34003, 22.46, 20.43269, 19.2456, 19.76627, 21.64799, 22.83505, 23.75811,
    24.08145, 21.84507, 20.51528, 25.59396, 28.70011, 26.54275, 31.31444,
    29.53227, 24.86761, 20.16363, 22.68626, 23.04077, 15.78924, 15.79892,
    15.25037, 15.09233, 14.05874, 13.62304, 13.3221, 12.6078, 12.50501,
    12.40103,
  21.42112, 20.85741, 18.17082, 17.40793, 18.09113, 18.85623, 19.79267,
    20.15373, 19.14544, 17.60932, 21.00746, 24.90881, 22.40626, 24.07229,
    28.13893, 26.34744, 24.44588, 22.22359, 24.85374, 23.51625, 18.19759,
    16.55916, 15.36504, 14.99065, 13.59401, 13.1768, 13.09514, 12.56846,
    12.4333, 12.34788,
  21.12238, 20.1891, 17.93633, 16.39754, 16.88592, 17.2057, 17.52916,
    17.50539, 16.73971, 19.08452, 23.14189, 21.21106, 18.92451, 20.50479,
    21.53754, 21.22087, 22.28816, 23.77443, 24.14088, 24.244, 22.12461,
    19.12086, 15.65971, 14.935, 13.91474, 13.15023, 12.89454, 12.59611,
    12.42826, 12.35702,
  19.8102, 19.52791, 17.7284, 16.17218, 16.21221, 16.49116, 16.45894,
    16.13741, 16.8865, 21.05866, 22.36647, 18.03493, 18.90228, 19.64771,
    19.02671, 18.51116, 18.99996, 19.82127, 19.93918, 20.90143, 21.94673,
    21.50489, 17.39347, 15.57557, 14.39184, 13.5309, 12.90976, 12.59537,
    12.43757, 12.36802,
  20.52962, 19.012, 17.52969, 16.55425, 16.48473, 15.89989, 15.90656,
    16.07673, 18.57935, 21.98816, 20.01317, 16.60431, 18.19909, 18.60851,
    18.02349, 17.46089, 17.09858, 16.87908, 17.53962, 17.93076, 19.5284,
    20.64013, 17.68021, 17.86603, 16.26687, 14.16664, 13.03981, 12.72448,
    12.45771, 12.36722,
  20.82829, 19.3404, 17.45692, 16.32725, 16.98196, 17.18955, 17.36486,
    17.19144, 19.6258, 21.26989, 17.73503, 16.24223, 17.18612, 17.50289,
    17.02368, 17.15693, 17.1778, 16.42375, 16.3041, 16.15425, 17.67353,
    18.36355, 15.61952, 17.85801, 18.14661, 15.21683, 13.20054, 13.23565,
    12.80725, 12.41201,
  20.64325, 19.4677, 18.26098, 17.74958, 18.38811, 18.6899, 20.33801,
    21.91586, 23.07501, 20.43573, 16.40816, 16.62829, 17.35014, 17.98443,
    17.70144, 17.79002, 18.23097, 17.33413, 15.97362, 15.95452, 16.79783,
    16.29388, 14.80709, 15.78885, 17.0734, 16.91022, 15.11656, 13.7594,
    13.29684, 12.61545,
  20.18785, 20.28582, 18.38048, 17.86004, 19.31464, 20.70443, 21.58405,
    22.48483, 23.69428, 20.84009, 16.1807, 16.89025, 17.70418, 18.46861,
    18.54087, 18.80978, 18.57964, 17.8035, 16.4789, 15.78315, 15.83262,
    15.42396, 15.40753, 15.10931, 14.78343, 16.55844, 16.76617, 14.81037,
    14.34146, 13.31025,
  20.49761, 21.967, 20.90878, 20.1974, 20.67212, 21.35518, 22.62115,
    23.73021, 22.34883, 19.76104, 16.59094, 17.37275, 18.47036, 18.7041,
    18.20951, 18.41397, 17.95946, 17.30638, 16.72702, 15.66462, 15.66128,
    15.87943, 15.19355, 14.30462, 13.9791, 15.08809, 16.80177, 15.99097,
    14.64803, 13.53704,
  21.89855, 23.42082, 22.44582, 21.09575, 20.78652, 20.39071, 23.54781,
    25.1549, 20.74256, 17.69541, 17.25544, 18.21545, 18.95468, 18.56877,
    17.86948, 17.61763, 17.13069, 16.82195, 16.47854, 15.42809, 15.63834,
    16.82429, 16.82374, 15.82999, 15.69392, 16.1006, 18.54145, 18.6346,
    14.78875, 12.75885,
  24.29592, 26.58048, 21.19123, 20.2798, 21.12578, 21.22177, 23.43295,
    23.15738, 18.16841, 16.80667, 17.44828, 18.27544, 18.4602, 18.04491,
    18.09203, 17.74367, 16.72241, 16.20837, 16.35962, 16.51376, 17.3027,
    18.14688, 17.80089, 17.03307, 16.87596, 17.24014, 18.39212, 20.60179,
    18.30036, 13.47578,
  22.77522, 21.68687, 20.7141, 24.91386, 25.13228, 24.08742, 24.26913,
    20.52212, 16.78617, 16.92222, 16.79423, 16.69312, 16.75793, 16.90956,
    17.63842, 17.84039, 17.45332, 17.49394, 17.21302, 16.92486, 17.43127,
    17.23379, 16.1071, 15.38977, 15.7234, 16.49109, 16.8908, 17.5927,
    17.96986, 14.64424,
  21.24537, 20.59611, 22.70742, 25.97158, 25.36817, 25.39768, 24.98073,
    19.98924, 16.41107, 17.08581, 17.2466, 17.63976, 18.21078, 18.40203,
    18.54118, 18.71595, 18.11455, 17.10977, 16.41817, 15.55834, 15.11671,
    14.96014, 14.57382, 14.30276, 14.61458, 15.41408, 15.90906, 15.16222,
    14.44766, 13.16813,
  16.58157, 16.65324, 16.69835, 16.73582, 16.70657, 16.69424, 16.70024,
    16.74077, 16.79701, 17.02608, 18.31745, 18.82594, 16.95382, 17.26574,
    17.59743, 16.95816, 16.79205, 16.86447, 16.93733, 17.61389, 18.29069,
    17.81827, 18.10378, 18.94373, 19.76418, 20.22864, 24.42761, 28.61032,
    21.63848, 18.73319,
  17.09098, 17.32673, 16.86703, 17.27002, 17.02719, 16.76438, 16.85576,
    16.9609, 17.13554, 17.54391, 18.40564, 19.37084, 19.78989, 18.86447,
    17.95783, 18.15024, 17.13878, 17.28553, 18.18789, 19.29057, 19.03108,
    17.91618, 18.47258, 21.13726, 28.14631, 33.09914, 29.83121, 36.96264,
    24.21016, 20.10483,
  17.09108, 17.13811, 16.98521, 17.06653, 16.86465, 16.77132, 16.85964,
    17.04864, 17.24781, 17.40902, 17.70289, 18.5104, 19.22908, 19.88137,
    20.0916, 18.35073, 18.11561, 18.98591, 18.96622, 19.31929, 20.68049,
    22.86252, 24.90753, 27.94021, 36.56867, 45.12519, 37.02362, 36.94875,
    23.70106, 21.34978,
  17.04708, 17.03498, 17.25445, 17.49842, 17.80489, 18.57899, 18.72887,
    18.26413, 18.31352, 19.02102, 19.64477, 19.90284, 19.60466, 19.03855,
    21.03896, 22.66205, 21.55565, 19.07778, 18.90509, 20.03789, 25.38319,
    30.01398, 28.26824, 36.06796, 44.36651, 39.44283, 45.259, 34.19916,
    23.42739, 19.57944,
  17.88365, 17.13679, 17.61338, 18.13759, 18.92748, 19.24776, 18.93526,
    18.85274, 20.13103, 21.75576, 21.41491, 20.1291, 19.3311, 20.0664,
    21.47633, 21.79898, 20.20148, 18.67778, 20.53876, 28.32893, 34.06171,
    26.80202, 27.32876, 31.4716, 34.18383, 34.29247, 33.62029, 36.55087,
    33.57546, 21.23035,
  17.53176, 17.59309, 19.19654, 21.23991, 21.17709, 19.85263, 19.61355,
    19.37222, 19.09035, 19.3965, 19.57027, 22.17837, 26.59911, 27.27925,
    29.99786, 35.75061, 41.1595, 35.7243, 28.10309, 32.3453, 30.13299,
    23.40007, 25.48636, 28.06844, 30.59606, 30.53788, 34.06958, 54.74445,
    49.32928, 20.64123,
  17.6628, 18.67784, 20.63385, 22.50314, 22.31517, 21.17103, 22.26613,
    25.89155, 27.33557, 28.13014, 29.06982, 28.52336, 26.56281, 27.18437,
    33.98768, 44.87125, 42.96346, 34.58889, 27.88681, 28.26356, 25.03188,
    23.21278, 25.08009, 30.30009, 34.6035, 32.75636, 42.86358, 63.80604,
    51.4285, 18.3998,
  17.99934, 19.37216, 21.57931, 23.36371, 22.57472, 25.36751, 31.43722,
    29.64102, 26.61777, 27.47817, 26.8972, 24.98699, 22.22424, 23.89935,
    28.90971, 33.34893, 31.01723, 29.06735, 24.45866, 24.22467, 22.9608,
    22.78529, 26.11943, 31.7854, 32.83599, 30.62003, 45.97047, 61.23078,
    33.58841, 18.79226,
  20.23534, 20.78915, 22.91825, 23.62714, 25.40749, 30.70917, 29.29269,
    25.84955, 26.50862, 26.34219, 24.45135, 21.49145, 21.47037, 29.66508,
    37.13747, 29.76227, 27.60255, 30.71426, 30.73573, 26.85696, 22.62346,
    26.32692, 34.87746, 38.1927, 31.10636, 35.18453, 47.74574, 45.77366,
    23.76433, 18.80284,
  24.33158, 28.8445, 31.40337, 34.49134, 36.39176, 33.29755, 21.97726,
    21.94574, 20.90421, 21.02352, 24.06158, 32.39892, 36.88015, 36.87872,
    32.35516, 32.04208, 34.09534, 35.3659, 32.76749, 28.25187, 28.74647,
    31.07417, 34.08526, 34.80933, 44.3339, 60.09344, 51.37854, 26.51773,
    19.56085, 17.10465,
  37.59639, 43.13789, 44.14354, 38.8605, 38.47326, 33.6795, 27.21451,
    30.6721, 34.73099, 41.29538, 49.18254, 35.26032, 30.08855, 28.95317,
    27.60022, 30.32827, 33.47225, 33.00053, 30.43726, 28.40992, 32.06494,
    33.14703, 28.86605, 26.42207, 33.88514, 40.55232, 30.58755, 18.32825,
    17.69885, 16.65804,
  57.25041, 44.56091, 43.98079, 43.77953, 42.82199, 34.76955, 42.48843,
    44.65295, 40.76217, 42.83146, 39.6989, 25.41559, 26.84939, 29.13168,
    28.7956, 30.94976, 30.38969, 29.58732, 28.26391, 29.62703, 33.22352,
    30.95621, 23.77215, 28.50637, 35.24429, 25.61504, 18.08957, 18.02377,
    17.85755, 17.02179,
  69.91106, 56.6345, 68.22734, 76.77008, 78.51988, 72.34664, 61.02171,
    45.33384, 47.04829, 36.94451, 28.50057, 24.13295, 31.94212, 36.7089,
    34.75692, 30.93827, 31.12461, 29.18628, 27.84853, 34.66694, 37.66177,
    27.17498, 24.0227, 31.21165, 36.25718, 21.62629, 17.67052, 18.41616,
    18.67027, 17.71278,
  77.53625, 89.65367, 91.87019, 94.33588, 87.55993, 80.21899, 72.12336,
    66.37753, 52.06624, 41.39576, 51.72914, 54.42208, 60.40107, 61.73484,
    53.8725, 40.50208, 32.44747, 35.20982, 38.86651, 41.21802, 35.3543,
    29.25532, 34.3937, 29.75786, 23.39253, 18.97783, 17.96469, 17.82565,
    18.31618, 17.77069,
  73.49364, 73.69469, 77.57021, 74.82851, 65.3409, 64.63359, 77.19522,
    75.62879, 63.19856, 67.1823, 70.76989, 60.77221, 54.56457, 59.73115,
    57.42042, 42.25581, 41.19925, 43.95145, 48.15266, 48.01274, 38.72207,
    36.80386, 32.1481, 22.84293, 18.23162, 18.61423, 18.04862, 17.60649,
    17.52932, 17.20288,
  67.37066, 66.75079, 65.74638, 59.26641, 55.76982, 60.97446, 76.80858,
    79.46447, 57.93962, 60.93998, 58.28716, 47.66686, 41.71724, 48.60915,
    45.65668, 42.56484, 46.32371, 43.5957, 42.71183, 43.05817, 32.13168,
    27.71709, 23.08168, 20.08616, 19.37659, 18.71502, 18.05988, 17.71171,
    17.34638, 16.96129,
  55.96358, 53.512, 47.82034, 45.4748, 45.33707, 48.45415, 54.55495,
    60.48929, 45.83974, 46.45892, 40.89923, 38.31338, 44.25009, 43.36034,
    42.33096, 43.21273, 43.69753, 38.98805, 38.91619, 38.51453, 23.95464,
    21.13187, 20.41724, 20.60123, 19.62573, 18.79771, 18.02101, 17.37946,
    17.16188, 16.93164,
  41.6838, 38.63638, 33.88774, 34.47335, 36.94935, 41.73073, 44.15583,
    43.48357, 38.25633, 34.45425, 34.63428, 42.9881, 47.08779, 47.42384,
    51.87198, 47.33352, 38.99393, 33.53489, 37.63858, 34.52943, 21.35643,
    21.95861, 21.54245, 20.91164, 18.7723, 18.29828, 17.98782, 17.042,
    16.92083, 16.79875,
  35.85873, 33.02151, 28.84637, 28.24524, 31.98717, 35.64897, 35.26134,
    32.16318, 28.94847, 27.95157, 35.37096, 42.11356, 38.85404, 42.55702,
    46.31256, 39.46251, 37.51863, 38.90166, 41.92456, 37.04469, 26.67786,
    24.85921, 22.40354, 20.69751, 18.17279, 17.79164, 17.65775, 16.98723,
    16.82795, 16.73485,
  33.39883, 31.68365, 27.9749, 25.44792, 28.38023, 29.54621, 27.39987,
    24.79517, 23.89732, 30.68416, 39.77935, 36.22163, 34.22657, 36.5671,
    35.79227, 31.66307, 33.4733, 38.72345, 40.82013, 40.35135, 35.20628,
    28.65687, 22.59109, 20.59335, 18.72462, 17.8085, 17.43718, 17.04171,
    16.81191, 16.74047,
  30.87923, 30.83896, 26.31335, 23.90576, 25.39098, 25.15143, 22.89344,
    22.16124, 25.35644, 34.54407, 37.67194, 30.85872, 33.13411, 32.37809,
    29.76175, 28.42922, 30.24697, 33.71922, 36.31073, 37.49681, 34.69343,
    30.59846, 25.02797, 21.53812, 19.30765, 18.3415, 17.4603, 17.05457,
    16.83644, 16.75934,
  31.27216, 29.45173, 25.66384, 23.97984, 23.96307, 21.57825, 21.25048,
    22.81656, 29.23287, 36.12323, 32.54794, 27.61313, 29.84027, 28.01573,
    26.16291, 26.58937, 28.48715, 30.85809, 32.79704, 32.39625, 30.39059,
    28.9171, 26.28812, 25.56203, 22.62754, 19.44374, 17.69177, 17.28854,
    16.88741, 16.77639,
  30.84233, 29.35321, 24.40135, 22.39786, 23.426, 23.60806, 24.36764,
    25.30027, 30.95841, 34.20713, 27.29433, 24.76103, 25.32352, 24.4128,
    23.89034, 25.9042, 28.78684, 29.40719, 29.10031, 27.59627, 26.89575,
    26.57313, 24.28493, 26.21532, 25.89467, 21.19366, 18.02589, 18.09733,
    17.39684, 16.85718,
  30.79472, 28.59983, 25.60402, 24.64475, 26.13619, 26.39268, 28.93151,
    30.8785, 34.23943, 32.16359, 23.84933, 23.41373, 24.00335, 24.82173,
    25.68369, 28.08742, 30.63071, 29.8779, 27.2967, 25.83771, 25.12848,
    24.22349, 23.25117, 24.23882, 25.1753, 24.172, 21.23373, 18.89571,
    18.03699, 17.13402,
  28.88823, 30.34507, 25.33573, 24.53492, 27.05055, 28.37904, 29.98213,
    31.67905, 35.6055, 31.76685, 22.09464, 23.08484, 24.70164, 26.73689,
    28.5234, 30.83637, 31.15418, 29.6621, 26.33117, 23.43374, 23.64616,
    24.00685, 23.48578, 22.24436, 21.27225, 22.98568, 22.96962, 20.27853,
    19.42974, 18.15014,
  30.72956, 33.64083, 29.61908, 28.16568, 28.99208, 29.46887, 31.32744,
    33.88382, 34.65032, 28.67389, 22.26783, 24.16259, 27.10555, 28.88769,
    29.20551, 30.28899, 29.5769, 27.71313, 24.94132, 22.06242, 23.61937,
    24.86806, 22.3955, 19.85366, 19.12239, 20.63617, 22.66189, 21.84727,
    19.73244, 18.36585,
  34.34735, 37.03201, 32.93685, 30.15916, 30.27685, 29.4316, 32.53349,
    34.27987, 30.72856, 24.68511, 23.55271, 26.48853, 29.08985, 29.47489,
    28.77379, 28.4129, 27.1806, 25.70341, 23.6975, 21.62722, 23.46773,
    25.73244, 24.41943, 21.93599, 21.29596, 22.1977, 25.19032, 25.33925,
    19.9816, 17.29881,
  37.94776, 39.84447, 31.96301, 30.08174, 32.66353, 32.53968, 34.45198,
    32.98343, 25.40608, 23.28371, 25.25494, 28.23966, 29.60826, 29.04763,
    28.68106, 27.53185, 25.42697, 24.15795, 23.31113, 23.27919, 26.1133,
    28.0506, 25.80409, 23.69864, 22.97146, 23.87406, 25.41681, 27.89716,
    24.8236, 18.41265,
  33.34323, 28.48088, 28.2028, 33.97123, 36.20467, 38.05075, 36.61757,
    29.12204, 22.91522, 24.48203, 25.55091, 26.49671, 26.8436, 26.69173,
    27.09752, 26.78712, 26.2212, 26.32917, 24.87053, 23.84299, 25.7366,
    25.44829, 22.84297, 21.37089, 21.70677, 22.9638, 23.66267, 24.20992,
    24.04351, 19.98889,
  29.64376, 28.03023, 31.61768, 34.60424, 34.05807, 37.01614, 38.13795,
    28.65418, 23.25982, 26.12726, 27.34072, 28.53809, 29.16639, 28.96391,
    28.40245, 28.32521, 27.42901, 25.55003, 23.53345, 21.83039, 21.54498,
    20.76629, 20.00933, 19.69028, 20.23873, 21.30918, 21.85011, 20.82329,
    19.53158, 17.81959,
  22.5086, 22.80147, 23.1109, 23.42822, 23.52543, 23.76434, 24.13635,
    24.68974, 25.42079, 26.67971, 29.12259, 29.21857, 24.94227, 26.096,
    26.54402, 25.24112, 25.56973, 27.01894, 28.93694, 32.17549, 34.34489,
    33.21566, 34.86811, 38.50678, 41.79041, 43.40472, 50.12468, 53.44968,
    33.09039, 26.43221,
  23.61907, 24.19526, 23.34802, 24.59241, 24.20015, 24.07021, 24.81397,
    25.48834, 26.35131, 27.48434, 29.26198, 31.47954, 32.47672, 29.78357,
    28.16819, 29.55766, 28.71423, 31.66575, 35.67897, 39.32796, 40.68204,
    41.77135, 45.43098, 53.87151, 62.10931, 59.25993, 53.63185, 57.2375,
    35.10036, 28.54431,
  20.87235, 21.04109, 21.33919, 21.77267, 22.02536, 22.5012, 23.00684,
    23.70341, 24.52179, 25.49752, 26.85461, 28.97249, 31.09154, 33.85264,
    35.99153, 34.75489, 38.05727, 42.96665, 47.05204, 53.10375, 61.53101,
    70.02407, 74.5742, 76.98213, 78.72435, 72.40824, 66.11478, 54.53616,
    35.28928, 30.74379,
  21.46576, 22.12346, 23.75076, 25.53437, 27.37761, 29.55502, 30.06878,
    29.92052, 31.24359, 33.1718, 33.94588, 34.56681, 35.83637, 37.62833,
    45.28303, 51.00806, 50.29102, 49.86527, 56.74342, 65.03304, 76.06145,
    79.62125, 76.27049, 83.91981, 83.96996, 80.57727, 71.97065, 52.33747,
    35.00373, 27.68056,
  25.55767, 24.89079, 27.51581, 29.28959, 30.77028, 30.62017, 30.50353,
    31.42697, 34.14906, 36.14952, 35.09948, 35.98929, 38.49095, 43.73462,
    49.92455, 54.70407, 55.14107, 53.2858, 60.13803, 70.46452, 73.36832,
    63.37218, 64.78167, 73.60664, 79.80922, 77.97854, 70.5836, 74.64845,
    64.08525, 36.19307,
  26.47965, 28.77956, 32.41593, 35.92832, 34.70173, 32.1585, 33.76319,
    35.77761, 38.40771, 44.07131, 52.48996, 66.28545, 80.23509, 81.19419,
    86.7749, 93.61002, 92.17833, 82.32052, 69.94669, 70.7271, 63.56981,
    55.98156, 63.56676, 71.63427, 80.18195, 80.24619, 77.25339, 91.29163,
    76.20898, 33.82697,
  29.4421, 33.79673, 39.1751, 45.12517, 48.77331, 53.81628, 64.19153,
    75.70308, 80.90309, 83.57365, 84.93818, 79.49768, 70.06522, 71.19456,
    73.18051, 75.62961, 74.67078, 65.89037, 56.80946, 58.44721, 56.49036,
    57.78065, 64.94867, 74.6901, 77.73488, 69.9514, 74.93938, 85.33348,
    64.13918, 25.72426,
  36.54023, 44.12585, 52.38368, 60.83969, 65.91325, 76.15272, 83.22115,
    69.43047, 59.77123, 59.8204, 54.75579, 48.85982, 44.0727, 45.3092,
    48.14056, 53.13155, 56.0155, 55.26493, 49.1749, 51.36498, 52.7602,
    57.25257, 66.11668, 73.04143, 69.42484, 65.82667, 77.286, 76.33864,
    50.63254, 26.77032,
  51.78405, 57.19835, 62.92186, 65.64238, 66.05635, 68.46052, 57.91131,
    51.56145, 52.82448, 52.1558, 49.85686, 49.21083, 53.44576, 67.24873,
    75.347, 59.90014, 62.08932, 70.06032, 71.48274, 64.73028, 62.40301,
    76.80499, 91.27635, 90.75884, 76.05899, 82.24913, 83.9453, 68.35574,
    35.59982, 26.74955,
  75.45487, 83.5582, 79.68758, 81.84575, 73.4848, 61.53677, 44.02725,
    52.54893, 56.36579, 66.69679, 79.12228, 91.99686, 91.21104, 86.01089,
    78.6934, 86.39792, 92.79796, 93.61887, 88.99356, 86.30049, 94.09811,
    95.53432, 91.25765, 80.12049, 85.36179, 95.99141, 78.85338, 43.69689,
    26.62666, 23.24585,
  94.94455, 89.63989, 88.24911, 78.43039, 89.64792, 91.12924, 89.37807,
    98.09538, 105.9962, 109.8821, 99.50121, 72.85323, 68.8378, 69.22639,
    72.45596, 80.10301, 86.34566, 86.96249, 84.9454, 85.77985, 96.62381,
    90.97813, 69.75861, 60.92208, 68.33641, 66.59654, 44.0494, 26.48322,
    25.16451, 22.92625,
  96.90651, 82.1871, 94.96584, 105.4344, 105.0108, 92.54056, 96.41301,
    90.83595, 81.14064, 68.24138, 59.8048, 54.57684, 61.84315, 68.78917,
    72.16656, 74.07166, 73.66296, 73.2481, 70.92735, 72.9454, 81.96036,
    74.50355, 56.63328, 66.13285, 68.18221, 46.05246, 25.82148, 27.73483,
    26.31255, 24.15907,
  121.9262, 123.1342, 126.9897, 128.4194, 127.569, 115.459, 91.85335,
    80.66652, 81.27873, 60.32592, 58.57529, 62.45656, 74.91462, 84.37593,
    81.46349, 69.8668, 71.60389, 68.31854, 66.47137, 73.3478, 76.7908,
    66.04276, 58.62156, 58.36454, 52.78847, 36.80207, 27.43301, 29.93811,
    28.87889, 26.03252,
  126.0984, 127.249, 126.4691, 124.0207, 114.374, 112.6086, 117.503,
    117.8905, 98.65152, 102.5441, 116.058, 111.5483, 120.3013, 121.8121,
    104.2433, 85.67319, 85.11679, 90.36749, 95.82073, 91.32394, 76.00353,
    61.59061, 56.1649, 43.33928, 34.87695, 31.39814, 28.32818, 27.43474,
    27.18469, 25.54697,
  107.0111, 97.38606, 95.51788, 95.12443, 98.7503, 110.5964, 121.6374,
    123.1659, 120.4775, 121.44, 120.5069, 114.8095, 119.1761, 120.3739,
    115.5353, 114.0894, 104.5829, 103.5352, 102.5064, 89.14282, 59.24047,
    52.85604, 40.94616, 33.63343, 30.96197, 29.78516, 27.6784, 26.03786,
    24.94878, 23.98068,
  90.31755, 91.07861, 94.95348, 99.27943, 104.1288, 115.8529, 123.7413,
    120.6722, 113.4384, 110.5769, 109.6263, 100.4899, 98.46533, 112.2028,
    109.6085, 105.9362, 103.2183, 88.98033, 78.0108, 64.21478, 42.17993,
    40.88837, 33.63786, 31.91086, 31.00128, 28.94184, 26.83267, 25.69567,
    24.49871, 23.6251,
  80.94949, 79.04677, 83.19867, 88.24945, 93.20025, 98.73604, 102.0869,
    102.0731, 97.57341, 95.0973, 89.04563, 100.371, 115.197, 107.2795,
    102.5443, 93.92816, 82.96629, 68.81773, 63.19765, 56.32303, 36.23933,
    37.96624, 33.97827, 31.80818, 30.416, 28.93717, 26.32748, 24.60371,
    24.05131, 23.59306,
  65.86634, 70.02328, 71.29402, 75.42169, 78.64786, 82.96976, 84.97808,
    85.62546, 87.01117, 86.97517, 101.8667, 120.7015, 121.3382, 117.0589,
    111.9765, 89.49342, 65.59074, 55.17142, 60.28162, 54.65193, 37.41383,
    38.89288, 35.02265, 32.97411, 29.20601, 27.55442, 26.13051, 23.76144,
    23.47257, 23.20344,
  73.67604, 72.1496, 63.47395, 60.23553, 63.12654, 65.65419, 69.48695,
    75.06155, 79.11054, 88.7656, 105.526, 107.0279, 90.28255, 90.19009,
    83.83809, 74.39494, 73.31326, 76.5081, 78.20206, 66.7106, 47.22182,
    40.8691, 35.67847, 32.38985, 27.94244, 26.23858, 25.32854, 23.68252,
    23.22247, 23.0847,
  70.36971, 64.69687, 54.5475, 48.25282, 51.70254, 56.06428, 62.77777,
    70.14976, 79.08275, 92.57478, 95.68411, 76.14098, 68.9482, 67.36341,
    64.05518, 64.63087, 71.18544, 78.65274, 78.05125, 71.71358, 58.07365,
    45.57613, 36.03253, 32.54988, 29.26014, 26.26399, 25.02312, 23.78707,
    23.17439, 23.11095,
  60.98682, 54.6631, 46.02228, 42.27735, 46.91312, 53.26602, 59.94091,
    66.77352, 74.59347, 80.65451, 71.78242, 55.9104, 61.09038, 61.61166,
    61.09766, 61.64947, 64.50748, 65.80229, 64.64131, 60.38728, 54.01077,
    50.28761, 42.55397, 36.01152, 31.54965, 27.73637, 24.99879, 23.87311,
    23.22529, 23.13825,
  58.41341, 48.89066, 43.94666, 43.62357, 48.52699, 51.42619, 57.67519,
    61.85845, 68.34357, 69.52567, 56.43289, 49.58899, 57.02745, 58.53897,
    57.89549, 57.45002, 55.49197, 53.05087, 51.45444, 49.29079, 48.39552,
    47.80585, 46.47392, 44.87622, 37.41044, 29.14762, 25.21523, 24.34951,
    23.32399, 23.14344,
  55.73632, 49.75963, 43.91237, 44.74757, 53.86979, 58.55502, 59.67794,
    57.56179, 59.59102, 56.67677, 44.75457, 47.52261, 52.64964, 54.55626,
    52.67691, 51.87292, 49.7417, 44.77985, 43.07536, 43.08791, 43.79428,
    43.76563, 42.3273, 43.0684, 41.48997, 32.76432, 26.83477, 26.51678,
    24.61781, 23.29857,
  58.67077, 56.31337, 56.15667, 60.09685, 65.40266, 66.35749, 68.16898,
    64.19833, 63.97185, 54.01228, 43.1041, 50.68041, 54.64201, 56.93908,
    54.56726, 52.55971, 51.08569, 46.67407, 42.40756, 42.26233, 42.00491,
    41.06599, 39.67884, 38.93325, 39.71122, 39.06469, 33.8399, 28.29316,
    26.32138, 24.03822,
  61.78323, 64.29487, 60.83762, 63.63778, 67.75071, 66.57008, 63.25724,
    62.88543, 66.81012, 56.7308, 44.93286, 53.37228, 57.03018, 58.7498,
    56.63382, 55.74479, 52.37524, 48.26526, 44.34291, 41.32294, 41.78305,
    41.96799, 39.48201, 36.5891, 36.12324, 39.73294, 39.83964, 33.51998,
    30.49701, 26.97864,
  73.62479, 79.06467, 77.10967, 71.69338, 67.43639, 64.23079, 68.20846,
    72.39701, 66.97856, 54.63083, 52.20058, 58.95546, 61.27554, 58.86219,
    54.17026, 53.14843, 51.27834, 48.60295, 46.22391, 42.84513, 42.73236,
    41.90416, 37.47953, 34.66045, 35.64737, 38.58384, 41.26416, 37.59647,
    30.33868, 26.68686,
  86.21266, 87.89532, 76.74583, 68.19363, 64.77573, 62.64672, 71.07626,
    71.58009, 59.84512, 52.67355, 57.67213, 60.62701, 59.98606, 55.96067,
    52.69138, 51.16209, 49.07972, 47.0497, 44.61455, 41.83776, 43.44822,
    46.82503, 46.26142, 43.47706, 43.52803, 45.43744, 49.07647, 45.37204,
    30.87355, 24.15575,
  89.61628, 83.27893, 71.70351, 71.15636, 72.31679, 71.92492, 73.1584,
    66.18655, 53.79071, 56.19123, 59.36157, 59.69081, 57.40631, 55.00615,
    53.67835, 50.61789, 46.70708, 45.59237, 47.35049, 50.37579, 53.64692,
    54.20213, 50.16805, 48.26274, 48.4936, 50.2913, 51.50761, 52.58103,
    43.63597, 27.71349,
  73.27715, 68.76983, 75.12307, 81.7612, 82.44965, 81.70877, 75.06802,
    58.74815, 51.35098, 53.7773, 50.17787, 47.97518, 48.19321, 49.78483,
    51.83334, 52.60915, 52.84778, 54.47748, 54.31728, 52.82118, 53.33,
    50.66512, 46.46365, 44.71587, 45.94367, 47.14069, 46.24029, 42.80302,
    38.92424, 30.87037,
  73.21827, 76.35086, 77.85464, 77.32137, 77.56264, 82.55293, 80.57944,
    61.12687, 50.25022, 53.73523, 54.98768, 58.8461, 62.21916, 63.01811,
    61.59269, 60.09181, 55.53659, 50.33201, 48.47998, 45.9416, 43.54,
    41.8299, 40.30693, 39.33228, 39.26869, 39.32133, 37.57333, 32.74307,
    28.40789, 24.33109,
  28.59611, 28.98289, 29.50935, 30.16899, 30.68094, 31.50916, 32.59768,
    33.90456, 35.48166, 37.59509, 40.51116, 41.51608, 39.45813, 41.27187,
    42.71281, 42.78656, 43.52652, 44.98155, 46.45382, 48.78421, 50.11272,
    48.97228, 50.10143, 52.6993, 54.2778, 53.73693, 57.71852, 58.50591,
    40.87623, 34.91395,
  29.23173, 30.03848, 30.07635, 31.89178, 32.55482, 33.71204, 35.90963,
    38.18796, 40.72073, 43.59586, 47.02406, 50.84816, 53.54743, 53.10834,
    53.34045, 54.83456, 54.2897, 56.02399, 58.10607, 60.18179, 60.72902,
    60.57547, 61.44981, 64.76685, 67.86544, 61.46291, 53.32217, 56.55197,
    41.67352, 36.44741,
  29.78407, 31.2143, 32.96396, 35.00518, 37.11072, 39.37751, 41.68129,
    44.21344, 46.86015, 49.44634, 52.12208, 55.29715, 58.3475, 61.59002,
    63.48893, 62.11953, 63.87822, 66.8, 69.58526, 74.32653, 81.46535,
    87.38126, 87.28289, 83.37654, 79.32169, 73.30316, 64.42974, 52.62915,
    40.32436, 37.21441,
  35.92013, 38.46434, 41.88543, 45.50887, 48.83707, 52.17439, 53.88963,
    54.91159, 56.79894, 58.38142, 59.15557, 60.08771, 60.5576, 60.7952,
    64.98758, 67.28964, 64.80236, 63.54929, 68.92487, 75.27719, 83.93944,
    85.17975, 80.52539, 85.67236, 83.82759, 81.58838, 76.30484, 59.76095,
    43.99026, 35.88128,
  42.71618, 45.19032, 49.73551, 53.64093, 56.84817, 58.82108, 60.60901,
    62.47634, 65.44135, 67.45027, 67.51165, 69.8525, 71.87476, 72.77131,
    73.90727, 74.44865, 71.4062, 67.12048, 69.44654, 76.06935, 76.37086,
    68.16507, 70.42556, 77.56793, 83.68582, 84.12305, 79.88343, 84.30999,
    73.66333, 45.22838,
  56.55286, 63.36744, 69.37181, 75.07704, 75.66794, 76.04111, 79.98778,
    81.47752, 81.86771, 84.53552, 89.99901, 100.3094, 109.9755, 106.7415,
    105.9732, 105.2328, 101.4176, 91.19679, 79.01559, 75.98371, 67.4362,
    60.54908, 66.63507, 71.82407, 77.19276, 76.7599, 75.7435, 88.72934,
    77.99358, 40.65639,
  68.44286, 74.61619, 79.62938, 84.6386, 85.99615, 88.1242, 94.91557,
    100.2808, 99.53247, 94.90372, 89.71115, 79.05098, 67.67386, 69.09353,
    70.13179, 71.85098, 72.7735, 68.9753, 62.97356, 63.69973, 61.93003,
    62.09401, 66.69962, 72.8311, 73.47565, 67.74769, 71.16185, 78.53375,
    63.7789, 33.09241,
  62.17052, 66.21661, 71.22439, 75.92694, 78.04369, 85.20995, 87.28413,
    70.53519, 63.10365, 64.7742, 62.99903, 61.85344, 61.4956, 64.38033,
    66.94901, 70.20968, 73.03909, 71.58691, 66.34491, 66.34576, 67.27641,
    70.81844, 75.9792, 77.98487, 73.74178, 72.81398, 79.01063, 74.23959,
    53.15977, 34.99452,
  69.96615, 73.03712, 76.68958, 79.25719, 81.97527, 85.16506, 77.10117,
    79.17588, 85.18947, 88.81799, 91.14467, 93.53609, 97.77001, 108.001,
    110.5945, 96.07894, 94.49874, 95.73395, 92.22516, 83.48969, 79.6358,
    87.15435, 94.5477, 90.27264, 79.43837, 83.85469, 80.92644, 64.26589,
    38.59715, 34.64573,
  99.67809, 106.961, 99.6814, 100.187, 101.7195, 96.12981, 80.30768,
    90.51468, 93.65406, 100.0779, 106.7332, 113.5504, 111.2956, 107.125,
    101.289, 105.2697, 105.5393, 101.6965, 96.80695, 94.39404, 95.18889,
    89.76341, 83.05035, 73.59568, 77.42887, 84.88599, 71.76186, 45.39617,
    34.01046, 31.97508,
  122.1322, 121.556, 119.8326, 108.2618, 116.2957, 111.9268, 104.9924,
    108.4323, 109.4165, 103.7092, 88.93031, 71.0474, 68.39121, 68.74808,
    68.77325, 70.23394, 72.98106, 73.45563, 74.10014, 78.22431, 87.17545,
    80.55783, 65.66589, 62.18016, 67.57936, 63.87564, 45.92195, 34.66679,
    34.45845, 32.13155,
  126.7541, 123.1424, 125.5411, 126.2118, 123.715, 103.2068, 101.6963,
    94.82175, 86.17004, 75.08461, 69.84789, 66.72779, 70.02965, 71.18398,
    67.97877, 65.53904, 63.3955, 63.69518, 64.67526, 69.68716, 78.33691,
    76.18483, 65.13214, 74.12408, 74.9704, 55.85952, 36.61477, 40.1922,
    36.18434, 33.65202,
  133.0197, 132.6437, 134.0821, 134.7417, 133.8158, 130.2484, 123.654,
    115.9198, 119.7935, 101.8069, 95.78098, 91.32124, 98.41838, 99.6664,
    86.56668, 70.99802, 71.6431, 69.28943, 68.02942, 71.93515, 73.32294,
    66.96477, 60.73088, 56.72386, 54.78783, 47.32797, 38.19806, 39.60093,
    38.60851, 35.20922,
  122.682, 123.2056, 123.4361, 123.392, 123.3848, 123.9935, 124.9044,
    125.3342, 123.8905, 124.4357, 125.2651, 123.6625, 124.924, 125.1335,
    112.9206, 90.59061, 85.12196, 87.5621, 88.3737, 79.57812, 65.93399,
    57.22425, 51.18676, 43.25241, 38.77403, 37.97155, 35.59622, 34.7206,
    35.23398, 34.30732,
  107.2776, 105.7406, 111.7342, 116.4781, 120.6503, 123.9044, 125.7634,
    125.5747, 122.8146, 121.2601, 111.6638, 102.8747, 103.5781, 103.7871,
    100.6838, 97.51505, 85.51059, 79.93504, 78.07399, 70.5528, 53.25903,
    52.12889, 44.33692, 40.91126, 39.39684, 37.39167, 35.74387, 34.28998,
    33.29525, 32.69683,
  105.645, 110.1327, 112.1234, 113.5304, 113.0571, 114.6181, 116.4461,
    108.1354, 96.86441, 91.30595, 88.58257, 80.85596, 77.01715, 84.23878,
    80.518, 76.88374, 76.61493, 67.68483, 63.45882, 57.34988, 45.40416,
    47.03265, 42.31525, 40.59424, 39.6254, 37.46367, 35.30251, 34.37993,
    33.47905, 32.71306,
  88.36859, 86.61529, 89.75186, 93.34132, 96.1978, 98.77576, 98.6599,
    97.01333, 92.85245, 87.228, 80.57881, 89.16507, 96.84173, 86.99342,
    80.37849, 73.25357, 67.6492, 62.74563, 62.45368, 58.24851, 45.49392,
    47.26298, 43.25509, 40.38941, 38.9206, 37.54107, 34.77598, 33.05124,
    32.9433, 32.60896,
  78.41968, 82.26186, 82.72135, 86.71484, 89.00566, 90.96162, 90.91422,
    89.83783, 90.58681, 89.28062, 99.00546, 107.6908, 104.0674, 100.2761,
    95.36922, 83.09982, 71.92665, 68.55748, 70.58851, 61.95277, 46.63162,
    45.75743, 42.72384, 40.83704, 37.33139, 35.89102, 34.89119, 32.52061,
    32.37571, 32.19535,
  91.74548, 85.4949, 73.91337, 67.59726, 68.30375, 67.13908, 67.99467,
    70.64616, 72.28329, 77.76568, 85.82748, 85.02976, 77.05814, 81.81164,
    84.09914, 86.52611, 93.85375, 98.50808, 92.52155, 79.02827, 58.30328,
    48.38624, 43.46429, 40.68908, 37.08658, 35.32666, 34.51702, 32.84228,
    32.33085, 32.21298,
  86.12501, 78.30099, 65.30981, 57.17122, 58.50806, 59.82832, 62.93949,
    66.27525, 71.21178, 78.11357, 77.71912, 66.41566, 66.14744, 65.70252,
    64.92349, 65.16494, 70.09007, 76.34758, 78.26247, 75.46992, 66.73632,
    56.38638, 47.3005, 43.6177, 40.05497, 36.11798, 34.55645, 33.0966,
    32.28875, 32.23121,
  77.38298, 69.00021, 58.15711, 52.8015, 54.76542, 57.24219, 59.64268,
    61.87124, 64.86367, 66.52541, 60.62635, 52.51678, 56.66586, 56.19698,
    54.46357, 52.91365, 54.29862, 57.07732, 60.32775, 61.96553, 62.59407,
    62.60399, 56.27378, 49.33897, 43.32486, 37.81092, 34.61618, 33.20341,
    32.3217, 32.25067,
  75.69099, 67.85014, 59.14315, 56.56446, 57.69336, 56.45705, 57.66451,
    57.55782, 59.99658, 59.34594, 49.94324, 45.98424, 49.21681, 49.19014,
    47.90213, 47.69987, 47.8092, 49.28032, 52.01748, 53.73709, 55.28126,
    56.36728, 57.63357, 56.34449, 49.09969, 39.79924, 35.50676, 34.23285,
    32.67542, 32.22421,
  78.21223, 74.63985, 66.19276, 62.75973, 66.74783, 65.57078, 62.22467,
    57.22316, 56.17329, 53.1233, 46.08941, 47.51729, 49.21375, 50.27732,
    49.00116, 49.76328, 49.81673, 48.11452, 48.73623, 49.8893, 50.89701,
    51.70731, 52.00595, 54.3989, 54.73682, 46.04912, 38.60735, 36.98315,
    34.56429, 32.43382,
  86.89266, 85.9234, 81.6105, 80.19772, 78.84977, 77.63101, 77.74268,
    74.16228, 73.73326, 65.72517, 58.02855, 62.17081, 64.06936, 65.95016,
    64.02913, 62.70996, 61.29782, 58.01969, 54.54885, 53.60037, 52.93835,
    52.35097, 51.94501, 51.65538, 53.42211, 53.65517, 47.20425, 39.94886,
    37.43405, 33.81232,
  84.77499, 83.0089, 74.52969, 73.0874, 74.09728, 72.28392, 71.93333,
    75.16359, 79.09572, 71.27335, 63.31495, 66.8851, 69.36463, 70.26519,
    68.4424, 67.43003, 64.18777, 61.78587, 59.66061, 57.08246, 55.83878,
    54.28588, 51.39181, 49.49002, 50.51052, 53.42019, 53.16227, 45.23332,
    40.17008, 36.2279,
  95.69542, 92.49114, 85.1498, 78.28897, 75.53046, 74.53276, 79.23325,
    81.94722, 77.4021, 69.93404, 68.68813, 70.8504, 72.00156, 70.53465,
    66.90023, 66.80042, 66.26234, 65.18103, 64.84652, 63.34333, 62.25338,
    60.50745, 56.09917, 52.82165, 52.96787, 53.83724, 54.5555, 47.7012,
    38.00259, 34.90202,
  97.24885, 91.45792, 81.44248, 74.75308, 72.74203, 69.53844, 74.97114,
    75.46517, 70.0845, 67.00895, 69.89009, 70.93183, 72.76788, 72.82012,
    71.64258, 70.99903, 70.03275, 69.86548, 70.16113, 70.28332, 70.95546,
    72.66809, 71.42706, 67.37417, 66.07735, 66.23157, 67.21296, 59.50541,
    41.96191, 33.06193,
  97.12329, 91.44958, 84.51401, 82.36205, 80.21839, 77.12721, 74.26923,
    69.78027, 63.9271, 66.65677, 69.18417, 72.71662, 73.99159, 74.81494,
    74.36907, 72.33572, 69.55721, 68.61877, 69.74878, 70.29227, 67.87636,
    64.12542, 60.56965, 59.72724, 60.36926, 61.44818, 62.30402, 62.99171,
    54.34142, 37.58578,
  81.77367, 80.21703, 83.1516, 84.84554, 86.73128, 86.4534, 79.61958,
    66.34248, 62.81641, 65.00858, 63.74408, 63.61362, 64.49206, 64.51795,
    64.23038, 62.96598, 59.61318, 56.91251, 53.57112, 50.37089, 49.49968,
    48.26889, 45.71063, 44.05038, 45.34068, 46.67312, 46.36655, 44.03102,
    43.62461, 38.9856,
  71.758, 73.38019, 72.97404, 73.03062, 78.05315, 85.52908, 84.52223,
    69.78334, 63.30535, 67.13622, 68.68613, 69.6031, 68.24803, 64.09753,
    58.89357, 54.63737, 47.57752, 42.04292, 41.20601, 40.36868, 38.90574,
    39.32805, 39.42392, 39.32542, 39.66634, 40.76747, 40.67619, 37.51897,
    34.33886, 32.19266,
  41.62434, 42.62966, 43.4259, 44.2993, 44.93496, 45.6127, 46.35691,
    47.08173, 47.84407, 48.87648, 50.35489, 50.4921, 48.53954, 49.05954,
    49.28967, 48.63865, 48.69717, 49.38861, 50.14616, 51.33061, 51.66921,
    50.41522, 50.93289, 53.02333, 54.62227, 53.76993, 55.5476, 56.37892,
    45.18091, 41.20069,
  47.05598, 48.35077, 48.61106, 49.98859, 50.32429, 50.92158, 52.04282,
    53.07924, 54.18075, 55.41512, 56.91625, 58.75417, 59.79593, 58.60653,
    57.85446, 58.17989, 57.52631, 58.59436, 59.88263, 60.86186, 60.96208,
    60.53857, 60.7939, 63.74794, 66.35063, 59.80909, 52.44327, 54.63987,
    45.48812, 42.01136,
  49.97999, 51.21634, 52.03248, 52.75125, 53.33585, 54.07652, 54.92669,
    55.93525, 57.02261, 58.0691, 59.20343, 60.69916, 62.10804, 63.76374,
    64.72038, 63.56509, 64.62465, 66.79121, 68.86051, 72.02711, 77.38441,
    82.1729, 82.15, 78.99942, 75.38498, 69.64759, 61.79853, 52.55189,
    44.68363, 42.67909,
  55.21225, 56.51378, 57.80535, 58.93107, 59.72408, 60.71348, 61.02407,
    61.06411, 61.76266, 62.39312, 62.43061, 62.53219, 62.33644, 62.06717,
    64.68392, 66.15192, 64.45592, 64.062, 67.86861, 72.23779, 79.04333,
    79.82561, 74.57825, 77.72728, 75.46213, 73.32648, 70.58322, 59.12494,
    47.74406, 42.11671,
  62.72818, 63.27891, 64.61996, 65.3083, 65.39423, 65.44503, 66.12886,
    66.54451, 67.9983, 69.07494, 69.2758, 70.74519, 71.53465, 71.07352,
    71.50396, 72.14716, 69.5042, 66.00573, 67.72142, 72.81383, 72.81847,
    64.92516, 65.96922, 70.92737, 75.38902, 76.3348, 75.31284, 80.88653,
    72.2173, 49.88632,
  69.18527, 71.86668, 74.20766, 76.21352, 75.25956, 75.04708, 77.67654,
    78.51057, 78.28583, 79.47791, 82.90273, 91.14045, 98.39738, 94.64256,
    94.64483, 95.0489, 91.03236, 83.4892, 74.72594, 72.55587, 65.24672,
    59.01331, 63.10244, 66.84381, 71.33904, 73.02251, 75.70825, 87.28429,
    77.06416, 45.7713,
  70.18172, 73.95406, 77.14931, 80.17235, 81.38968, 84.32392, 91.06802,
    96.55904, 96.03246, 91.48444, 86.43223, 76.93507, 66.84246, 67.07898,
    67.82989, 69.37207, 69.82944, 66.54767, 62.92, 63.33939, 61.39109,
    60.36958, 63.03853, 66.92874, 67.61657, 65.28479, 70.07214, 77.28763,
    64.07691, 39.82464,
  74.86263, 79.16626, 82.68421, 85.67017, 86.82404, 91.87331, 93.86053,
    80.85413, 73.80363, 73.49275, 70.19615, 67.20638, 65.10467, 65.13947,
    65.49551, 67.04779, 68.83384, 67.66211, 64.45465, 64.43309, 64.63827,
    66.4855, 69.56629, 71.13542, 68.90785, 69.56837, 75.6703, 72.96191,
    55.48653, 40.90308,
  86.74518, 88.80152, 90.15916, 90.84782, 91.86642, 91.82581, 82.45605,
    81.93396, 84.23318, 83.77071, 82.91472, 81.99702, 82.3758, 87.72938,
    89.0062, 80.41515, 79.95439, 81.10634, 79.03111, 73.9729, 71.21954,
    75.36394, 80.32292, 78.30118, 72.4854, 77.17721, 77.90051, 64.49553,
    43.62689, 41.07994,
  98.39018, 100.3571, 94.60281, 93.99951, 94.28184, 87.26581, 71.52849,
    77.08547, 76.52238, 78.3726, 80.386, 83.39831, 82.587, 80.87941,
    78.60409, 82.28957, 83.41023, 82.52785, 81.05893, 81.01784, 81.49017,
    77.56326, 72.9631, 67.07666, 71.39805, 79.38756, 70.32549, 49.69181,
    40.6645, 39.34302,
  119.629, 118.8925, 113.4661, 101.1488, 102.8734, 93.07621, 84.08456,
    84.78662, 85.60193, 81.50102, 70.84924, 59.80345, 58.49712, 59.73448,
    60.7369, 62.33824, 64.77652, 66.35898, 68.18721, 71.83214, 78.05103,
    74.21721, 64.0219, 62.36866, 66.65524, 64.27639, 50.39421, 41.25532,
    41.16224, 39.48088,
  126.8893, 124.2346, 125.5834, 124.7136, 121.6341, 98.69383, 92.96745,
    84.57889, 78.02299, 71.49409, 66.71039, 63.9495, 65.96674, 65.81084,
    62.26804, 61.11692, 60.17675, 60.57709, 61.89976, 65.78757, 72.08115,
    70.5594, 63.46293, 69.89845, 71.4426, 57.27118, 42.93594, 45.29623,
    42.3463, 40.46965,
  129.9945, 130.35, 131.0573, 129.8775, 127.3938, 123.692, 117.5527,
    105.4982, 106.894, 94.36238, 87.59997, 82.67919, 87.37723, 88.44258,
    78.10739, 65.5229, 66.49668, 65.52815, 64.64779, 66.79195, 67.99828,
    64.64613, 60.29282, 56.68354, 55.26714, 50.24844, 43.88153, 44.74424,
    44.01886, 41.60206,
  119.5789, 120.3639, 116.27, 113.2715, 111.6302, 117.8223, 118.8991,
    117.6669, 107.8721, 108.9639, 111.7352, 106.3516, 105.7937, 104.9793,
    94.67759, 80.35312, 74.59138, 78.64473, 80.49109, 73.89207, 64.76155,
    58.65905, 53.62221, 47.15413, 43.55188, 43.35742, 41.97414, 41.31108,
    41.60847, 40.85031,
  85.17961, 81.29251, 82.92053, 83.27113, 84.9929, 88.87577, 94.44519,
    92.39703, 88.02924, 87.34219, 83.69817, 79.87273, 82.34026, 85.67374,
    84.9389, 82.59921, 76.29199, 72.60526, 72.12193, 67.52573, 56.13287,
    53.77038, 47.89012, 45.04552, 44.41716, 43.35069, 42.03868, 40.8961,
    40.15991, 39.77843,
  81.26019, 83.10104, 83.30222, 82.96777, 82.16714, 83.52068, 85.92065,
    82.53085, 77.04208, 74.0973, 72.48771, 69.33399, 68.37109, 72.60036,
    70.31915, 69.05551, 69.43049, 63.95065, 61.1142, 56.53815, 49.2652,
    49.53064, 45.88374, 44.70319, 44.39579, 43.31271, 41.80388, 40.91709,
    40.26593, 39.75345,
  72.92699, 71.73293, 72.82858, 74.60042, 76.18903, 77.55843, 79.78876,
    81.8956, 80.343, 76.6451, 72.17715, 77.74113, 83.12817, 78.00554,
    71.91276, 67.46626, 63.3759, 60.74627, 60.00396, 56.3219, 48.7422,
    49.35779, 46.47202, 44.49444, 43.81033, 43.18768, 41.34235, 40.04577,
    39.90294, 39.67928,
  68.42322, 69.3558, 68.44996, 70.37065, 72.31483, 75.09285, 77.22215,
    79.15122, 80.52031, 79.62853, 84.77866, 89.39271, 87.83609, 86.47669,
    83.0204, 76.2084, 70.5858, 68.6246, 68.09362, 61.02018, 50.36233,
    48.46753, 46.32225, 45.10388, 43.02003, 42.17, 41.29878, 39.69689,
    39.52284, 39.40152,
  75.95448, 70.58939, 62.4563, 59.06066, 61.47759, 62.46239, 64.13998,
    65.8343, 66.35233, 68.9951, 73.27472, 72.25357, 67.93944, 70.63757,
    71.8895, 75.01299, 81.29877, 85.51048, 82.85179, 73.21589, 59.23001,
    51.0077, 47.10144, 45.49599, 43.18803, 41.87206, 41.15282, 39.92512,
    39.50341, 39.44828,
  68.62766, 63.53449, 55.42895, 51.22099, 52.84791, 53.9233, 55.27953,
    56.74682, 59.46459, 63.88161, 63.92114, 58.35236, 58.82943, 58.15181,
    57.62853, 58.34729, 62.58421, 67.92655, 69.53165, 68.29549, 62.9229,
    55.92281, 49.82818, 47.30795, 45.04754, 42.52641, 41.29598, 40.08003,
    39.49965, 39.46312,
  63.68521, 58.95049, 51.16826, 47.41495, 48.42489, 49.41814, 50.7458,
    52.41345, 55.01031, 57.38261, 54.9313, 51.8999, 55.06772, 54.77351,
    53.49177, 53.15723, 54.66064, 56.97575, 58.85239, 58.96165, 59.12235,
    59.03931, 55.18076, 51.15704, 47.33262, 43.67037, 41.2781, 40.19217,
    39.54716, 39.47385,
  66.53957, 62.66905, 55.30422, 52.31933, 52.62302, 51.52355, 52.35505,
    53.13937, 56.08268, 56.6305, 51.84887, 49.95033, 52.03863, 52.11026,
    51.51718, 51.81984, 52.02414, 52.87516, 54.44164, 55.13607, 55.16989,
    55.00763, 55.49845, 54.72547, 50.79533, 44.89545, 41.9304, 40.87303,
    39.79064, 39.48729,
  74.12991, 73.71076, 66.02232, 63.36121, 65.34478, 64.97367, 63.11127,
    60.57352, 60.76165, 58.9098, 54.53133, 55.27195, 56.20387, 56.26456,
    55.09964, 55.41183, 55.143, 53.65703, 53.63754, 53.69854, 53.29953,
    52.67809, 52.29142, 53.75532, 54.33519, 49.10664, 44.18887, 42.77475,
    41.05251, 39.62427,
  80.33499, 80.39196, 76.69469, 75.67587, 75.58374, 73.69771, 73.97845,
    73.58614, 74.82767, 69.86016, 65.05182, 67.28661, 68.57513, 68.67061,
    66.68156, 65.11593, 63.51355, 61.05722, 58.38458, 56.61857, 54.75951,
    53.39434, 52.60843, 52.38125, 53.77921, 54.23747, 49.95008, 44.88974,
    43.04736, 40.51366,
  81.35023, 78.3061, 72.62575, 71.27293, 71.40958, 70.10426, 71.29331,
    75.3619, 79.23595, 74.00086, 68.07652, 70.19501, 71.47963, 71.62569,
    70.31379, 69.04902, 66.20721, 63.92866, 61.89532, 59.2799, 57.40689,
    55.06157, 52.36722, 50.72741, 51.67341, 54.07989, 53.93388, 48.21016,
    44.78758, 41.9953,
  87.37728, 85.24402, 80.30015, 75.44891, 72.85958, 72.04837, 76.30269,
    80.64527, 79.51347, 74.24107, 73.18379, 73.81303, 74.49097, 73.15589,
    70.9798, 69.90108, 68.17103, 66.76099, 65.98363, 64.07423, 62.57432,
    60.28131, 56.32162, 53.52359, 53.64659, 54.43486, 54.6879, 49.59647,
    43.19112, 41.14744,
  90.02831, 86.62515, 79.10429, 74.44904, 71.52715, 69.04082, 72.73928,
    74.25024, 71.74908, 69.60692, 70.91215, 71.72762, 72.13571, 71.93414,
    70.94495, 69.57747, 67.99091, 67.77835, 67.81967, 66.99226, 66.27369,
    66.41022, 64.88189, 62.13645, 61.43985, 61.82069, 62.45269, 56.93167,
    45.57893, 40.0261,
  84.58197, 82.38194, 78.09148, 75.76741, 74.35367, 70.09708, 67.79454,
    64.43358, 60.00281, 60.63779, 61.50494, 62.91385, 64.3933, 65.24983,
    65.58738, 64.7216, 63.16694, 63.32964, 64.86996, 65.19972, 63.13004,
    60.17602, 57.79049, 57.18634, 57.92841, 58.61678, 58.83445, 59.4898,
    53.67414, 42.89067,
  67.13869, 66.75912, 68.39249, 69.27161, 71.0599, 71.69331, 65.18055,
    56.0667, 53.0553, 54.13125, 53.64853, 54.07901, 55.11248, 55.75522,
    56.13174, 56.11969, 54.90079, 54.56246, 53.62246, 51.91718, 51.45121,
    50.65377, 48.96181, 47.93234, 48.6935, 49.17937, 48.57871, 47.24936,
    47.15644, 43.84195,
  55.88862, 56.39684, 56.00392, 55.24043, 57.87996, 62.90646, 62.46939,
    53.74242, 50.03701, 52.88618, 54.83636, 56.54046, 57.09528, 55.50531,
    53.2962, 51.40476, 48.09554, 45.36372, 45.32104, 44.88708, 43.99032,
    44.38836, 44.69398, 44.70701, 44.80696, 45.23949, 44.89959, 43.16544,
    41.23244, 39.55426,
  45.29335, 45.58469, 45.89895, 46.26022, 46.55883, 46.85506, 47.11548,
    47.41465, 47.83199, 48.61631, 49.89386, 49.73207, 47.66082, 48.28112,
    48.66629, 48.30045, 48.57813, 49.40085, 50.41115, 51.76444, 52.17982,
    51.19826, 51.78915, 53.63276, 55.20998, 55.16413, 57.04356, 57.8713,
    49.50937, 46.20861,
  48.89574, 49.33349, 49.09565, 49.81649, 49.77798, 49.84712, 50.1629,
    50.40674, 50.75249, 51.32278, 52.21123, 53.19686, 53.64138, 52.61024,
    52.22433, 52.8643, 52.5713, 53.8028, 55.32343, 56.50749, 56.83136,
    56.90961, 58.22092, 61.58344, 64.4867, 60.19243, 54.02582, 56.81538,
    49.51127, 46.77312,
  51.56903, 52.04779, 52.35212, 52.71784, 53.10713, 53.59303, 54.00613,
    54.57009, 55.22313, 55.88302, 56.73759, 58.02039, 59.31512, 60.95707,
    61.98788, 61.38914, 62.5438, 64.62553, 66.55956, 69.47046, 74.50359,
    79.58592, 80.08434, 76.437, 72.95335, 68.41669, 62.37384, 55.72668,
    49.34766, 47.63701,
  55.63955, 56.47929, 57.52077, 58.59272, 59.53217, 60.62953, 60.92953,
    60.90065, 61.50617, 62.22192, 62.64365, 63.62155, 64.1004, 64.15068,
    66.7933, 68.14249, 66.71942, 66.70242, 70.00029, 73.91297, 79.92548,
    79.86073, 73.88321, 75.39682, 72.11655, 70.47005, 69.30855, 59.43552,
    50.45518, 46.78645,
  58.44899, 58.50761, 59.61288, 60.46199, 60.95591, 61.26163, 61.84203,
    62.34455, 63.63025, 64.34938, 64.38747, 65.741, 67.05972, 67.92743,
    69.22058, 70.54037, 69.67963, 68.55905, 71.25307, 76.12341, 75.93592,
    67.93983, 67.55058, 71.44718, 74.47379, 75.04756, 74.07361, 79.03607,
    74.1721, 54.88,
  64.66405, 66.96911, 69.41421, 71.65829, 71.68687, 72.52888, 75.54935,
    77.05817, 78.33928, 80.82248, 84.98106, 94.07042, 101.967, 98.89308,
    98.94276, 99.25452, 95.74003, 89.03913, 81.45061, 78.09611, 70.67101,
    64.33784, 68.08289, 70.883, 74.63679, 75.80968, 77.19705, 87.84753,
    80.93742, 51.37631,
  71.97887, 75.24015, 78.19661, 81.10741, 82.54497, 86.07645, 93.43309,
    99.45459, 99.49208, 95.56055, 91.13786, 82.83693, 73.60487, 73.74838,
    74.45431, 75.40413, 75.47914, 72.2636, 67.73872, 66.68052, 63.96857,
    63.0931, 65.85992, 69.45989, 70.68318, 69.49772, 73.88943, 80.60876,
    68.40294, 45.07027,
  70.76889, 73.30738, 75.85839, 78.2135, 79.14232, 83.80134, 85.90269,
    73.6192, 66.61702, 66.20513, 63.32053, 60.85269, 59.56205, 60.48227,
    61.89051, 64.36887, 66.77405, 66.25321, 63.56095, 63.36124, 63.53528,
    65.22765, 68.45117, 70.85138, 70.4004, 72.26193, 79.23648, 77.29506,
    60.06575, 45.65114,
  75.00959, 76.601, 78.19522, 79.2755, 80.99255, 81.36024, 72.83578,
    71.63466, 73.62895, 73.41729, 73.34802, 73.49065, 75.00445, 80.07249,
    81.86301, 75.85655, 76.56087, 78.49141, 77.10175, 73.08785, 71.29091,
    75.13286, 79.26782, 77.57621, 73.71024, 78.78917, 80.41759, 68.9119,
    48.58778, 46.18559,
  86.01641, 89.79197, 86.58577, 88.22146, 90.94309, 85.08474, 71.2664,
    77.0041, 77.23492, 79.47419, 82.07135, 85.99994, 85.80527, 84.1768,
    81.59244, 83.97951, 84.74895, 83.43731, 81.73048, 81.01092, 81.43877,
    79.15291, 76.14223, 71.37866, 75.63167, 83.0248, 74.75472, 54.35633,
    45.64294, 44.82241,
  108.344, 106.672, 103.3571, 94.47404, 97.5583, 89.48114, 81.07023,
    83.97651, 84.7755, 82.29992, 74.43443, 65.18512, 64.51177, 65.39396,
    65.42773, 66.72723, 68.41214, 69.03678, 69.87301, 72.28746, 76.64215,
    73.59011, 66.33929, 65.38094, 70.40023, 69.10151, 55.25051, 45.70147,
    46.15784, 44.81578,
  112.826, 109.9119, 111.5271, 111.7877, 105.1801, 87.03619, 84.54634,
    78.00548, 72.22408, 68.59707, 64.91729, 63.45207, 65.61288, 65.61475,
    63.70665, 63.13208, 62.64196, 63.28111, 64.38002, 67.27589, 72.45679,
    71.77045, 67.01663, 73.11848, 74.26762, 60.52224, 46.86894, 48.93106,
    46.70292, 45.46983,
  119.4079, 119.3235, 120.1191, 119.4764, 117.6157, 113.8693, 103.2574,
    89.80712, 94.39681, 83.76595, 78.79889, 76.06185, 81.019, 82.24264,
    74.66207, 64.61418, 66.35141, 66.21026, 66.44238, 68.98674, 71.36295,
    69.77235, 66.62389, 63.97919, 61.39059, 55.03906, 48.26456, 49.09032,
    48.14938, 46.39132,
  111.6194, 111.422, 110.7019, 108.9421, 107.6342, 107.5345, 107.7369,
    107.0997, 101.5244, 101.3456, 105.6369, 102.3432, 100.5406, 100.7979,
    91.18564, 79.31741, 75.03264, 79.3531, 81.0787, 74.85725, 67.566,
    62.94052, 59.09802, 52.82281, 49.21325, 48.75825, 47.46593, 46.73681,
    46.75266, 46.04362,
  88.56085, 84.77819, 86.44363, 86.45119, 87.72395, 90.81933, 95.66444,
    94.61131, 90.27243, 90.11368, 86.75031, 82.92831, 84.67128, 86.39583,
    85.97207, 84.13082, 78.33725, 74.95947, 73.63461, 68.95447, 59.15336,
    56.89282, 51.79542, 49.41441, 48.98892, 48.29668, 47.2484, 46.18457,
    45.52438, 45.14652,
  78.6898, 80.62397, 81.3429, 80.68413, 79.70128, 80.88615, 82.65344,
    80.53649, 76.33934, 73.65452, 72.97987, 70.69029, 69.89583, 73.70037,
    71.97164, 70.85538, 71.00307, 66.28704, 63.65169, 59.16888, 53.00915,
    53.09937, 50.04346, 48.8598, 48.75321, 48.17604, 47.10524, 46.25554,
    45.60741, 45.13422,
  69.52666, 68.43285, 69.084, 70.13255, 71.29337, 72.35844, 74.01286,
    75.8522, 74.72597, 71.9521, 68.47195, 72.58676, 77.22596, 73.7778,
    69.74864, 67.04628, 64.43475, 62.31264, 61.58758, 59.05893, 52.87832,
    53.10697, 50.3373, 48.80813, 48.57501, 48.21727, 46.75336, 45.57621,
    45.3069, 45.05766,
  66.45657, 67.28698, 66.58906, 67.83144, 69.12727, 70.882, 72.32819,
    74.08306, 74.88647, 73.98486, 77.50121, 80.59369, 79.41427, 78.34325,
    74.13471, 69.1666, 64.9287, 64.18772, 64.70604, 60.53232, 53.10868,
    52.16485, 50.38305, 49.39354, 48.05179, 47.30489, 46.47748, 45.14249,
    44.97678, 44.84918,
  75.36086, 71.07139, 64.3192, 61.37608, 63.31236, 64.01989, 65.47562,
    66.87692, 67.24241, 69.44413, 73.04945, 72.13523, 68.07623, 69.7383,
    70.54028, 72.81218, 77.97842, 81.9058, 79.61285, 71.7326, 60.58361,
    53.999, 51.0645, 49.9744, 48.1181, 47.05027, 46.31609, 45.2581, 44.94611,
    44.86483,
  71.95602, 67.85081, 61.50118, 57.96555, 59.814, 60.83711, 62.16645,
    63.47908, 65.50589, 69.10619, 69.59552, 65.38988, 65.57655, 64.9229,
    64.18967, 64.49153, 67.47147, 71.42265, 71.89088, 69.17075, 63.40556,
    57.45395, 52.99431, 51.45359, 49.72236, 47.65832, 46.5456, 45.43306,
    44.93464, 44.90559,
  67.93914, 64.51984, 57.91836, 54.68325, 55.74747, 56.45963, 57.48969,
    58.65448, 60.51877, 62.53042, 60.65842, 58.07121, 60.62618, 60.50629,
    59.31583, 58.88781, 59.94256, 61.357, 62.15004, 61.18317, 60.35831,
    59.7875, 56.88709, 54.06395, 51.25031, 48.41562, 46.53773, 45.55162,
    44.96727, 44.89524,
  66.5679, 63.44967, 57.38839, 54.70572, 55.07563, 54.17535, 55.01414,
    55.71677, 57.98997, 58.59029, 55.04407, 53.42118, 55.30222, 55.65701,
    55.55254, 56.11149, 56.56131, 57.1236, 57.97501, 58.14291, 58.01694,
    57.74027, 57.67014, 56.72234, 53.37943, 49.05194, 46.89342, 45.94413,
    45.12482, 44.90376,
  69.34189, 68.55104, 61.38545, 59.03452, 60.66669, 60.44538, 59.11894,
    57.18709, 57.58192, 56.42582, 53.21087, 53.90593, 54.99517, 55.6149,
    55.51139, 56.48923, 56.90535, 56.04998, 56.02433, 56.01379, 55.77552,
    55.26117, 54.64441, 55.40667, 55.56445, 51.54434, 48.20044, 47.32101,
    46.00588, 44.97712,
  76.49056, 76.52067, 71.97247, 70.22449, 70.15181, 68.81738, 68.71446,
    68.09039, 69.30972, 66.1321, 62.62643, 64.51369, 65.83604, 66.28319,
    65.29707, 64.47914, 63.41677, 61.33923, 59.1539, 57.75354, 56.34929,
    55.5717, 54.74459, 54.38384, 55.26543, 55.03225, 51.80476, 48.47628,
    47.27268, 45.59488,
  78.72378, 75.16335, 69.71972, 67.5918, 67.68674, 66.87695, 67.74718,
    70.92774, 74.2657, 70.09586, 65.77688, 67.912, 69.23322, 69.86181,
    69.18533, 68.59283, 66.8007, 65.11781, 62.95852, 60.56804, 59.27688,
    57.75735, 55.49697, 54.07921, 54.68364, 56.00543, 55.39057, 51.35658,
    49.05109, 46.91553,
  83.57497, 80.44461, 75.1918, 70.41562, 68.70024, 68.27885, 71.74574,
    75.65062, 74.66376, 69.79652, 69.22967, 70.45806, 71.38883, 70.6996,
    69.15729, 68.45542, 67.78915, 66.78433, 65.1219, 62.87003, 61.71487,
    60.10076, 56.51458, 54.48133, 54.56956, 54.84657, 55.29765, 52.42987,
    48.13859, 46.2965,
  84.99175, 81.00498, 75.52986, 71.71846, 70.10666, 68.88499, 72.37025,
    73.85555, 72.16908, 70.11519, 71.26863, 72.103, 72.60658, 72.31995,
    70.97167, 69.87672, 69.21787, 68.94803, 67.64178, 66.29071, 66.6879,
    67.05038, 64.62497, 61.3386, 59.93685, 59.90427, 60.48982, 57.25136,
    49.33784, 45.30167,
  80.56327, 78.76997, 76.21417, 75.4701, 75.69825, 74.2478, 73.59612,
    71.49255, 68.75241, 69.4872, 70.55862, 71.79709, 73.0153, 73.59095,
    73.05004, 71.69152, 70.69559, 70.16862, 69.66042, 69.26899, 68.17855,
    66.05141, 62.6876, 60.84702, 60.29689, 60.35464, 60.47771, 60.71213,
    56.09635, 47.51108,
  67.72672, 68.16904, 69.38514, 70.45599, 72.46288, 74.36283, 70.51755,
    63.56468, 61.44653, 62.38181, 62.20554, 62.71976, 63.92629, 64.96873,
    65.39249, 65.33686, 64.65266, 63.99229, 61.93482, 59.78888, 58.85751,
    57.4968, 55.64737, 54.38351, 54.45522, 54.3227, 53.3998, 52.20569,
    51.69871, 48.4806,
  62.50801, 63.11036, 63.22066, 62.96919, 65.35766, 70.1225, 70.39114,
    63.15315, 60.03698, 62.25649, 63.85941, 65.26304, 65.24616, 63.54065,
    61.21733, 59.38021, 56.39747, 54.09177, 53.85361, 52.88239, 51.74132,
    51.77942, 51.72453, 51.44884, 51.12811, 50.71328, 49.68008, 48.19519,
    46.68399, 45.0832,
  38.54531, 38.58191, 38.65922, 38.79045, 38.90043, 38.96102, 39.10407,
    39.40165, 39.77732, 40.36547, 41.31208, 41.08038, 39.46223, 39.85838,
    39.99045, 39.44522, 39.37561, 39.57872, 39.89213, 40.64437, 41.04939,
    40.45446, 40.78252, 42.25909, 43.90136, 44.33519, 46.13856, 47.57794,
    41.8777, 39.38195,
  40.34765, 40.55698, 40.25793, 40.75923, 40.66934, 40.58554, 40.92001,
    41.29769, 41.72623, 42.23288, 42.75295, 43.1607, 43.24849, 42.29622,
    41.71379, 41.84103, 40.93742, 41.33812, 42.08205, 42.84266, 43.21305,
    43.83989, 46.01122, 50.70105, 54.80359, 51.01953, 45.30921, 47.965,
    42.22045, 39.94244,
  41.51162, 41.6292, 41.66489, 41.78375, 41.88912, 42.07094, 42.3284,
    42.70754, 43.13544, 43.54887, 43.95521, 44.56455, 45.13331, 46.05051,
    46.68695, 45.9678, 46.5645, 48.0196, 49.62383, 52.59199, 57.93347,
    64.34183, 67.00588, 65.67213, 63.34384, 57.85305, 52.58016, 47.27771,
    42.18621, 40.69212,
  44.52509, 45.2468, 46.18948, 47.13745, 47.89867, 48.80931, 49.0987,
    49.10558, 49.65914, 50.3351, 50.69027, 51.4925, 51.99838, 52.34219,
    54.75589, 56.21603, 55.41454, 55.68833, 59.16547, 63.84886, 70.53918,
    70.78082, 64.74927, 65.24004, 61.52031, 59.53829, 58.49372, 49.74146,
    42.21439, 39.68636,
  49.81944, 50.3098, 51.45898, 52.17965, 52.29605, 52.21253, 52.28021,
    52.11632, 52.62503, 52.66648, 52.35659, 53.56835, 54.97914, 56.38645,
    58.13839, 59.89645, 59.75876, 59.2441, 62.36524, 67.43924, 66.98383,
    57.81699, 55.49638, 58.87332, 60.95215, 61.21341, 61.25816, 66.62401,
    63.74156, 47.44119,
  52.17091, 53.18555, 54.51114, 55.52087, 54.60806, 54.40639, 56.50014,
    58.11604, 60.3517, 64.04498, 69.68224, 80.42366, 89.66645, 86.93965,
    87.42297, 88.68835, 85.19821, 78.53526, 71.61098, 68.24864, 60.53523,
    53.42776, 57.6321, 61.05869, 65.09249, 66.75987, 69.00569, 79.12297,
    72.56158, 44.93849,
  57.32599, 60.24128, 63.39376, 66.86481, 69.81821, 75.6786, 86.11546,
    95.88261, 97.87168, 97.39831, 96.89325, 92.70702, 83.32094, 82.07486,
    81.22706, 79.86053, 77.3356, 70.48457, 63.73244, 61.50761, 57.70966,
    56.8191, 60.07432, 63.61776, 65.18465, 64.52526, 68.74101, 74.53872,
    61.07281, 38.47498,
  69.38786, 74.72993, 79.67451, 84.98033, 89.06923, 96.92878, 99.84679,
    91.11156, 83.13484, 80.26077, 74.41003, 68.42978, 64.19092, 63.08952,
    62.48352, 63.15421, 63.1752, 60.52151, 57.34322, 56.72565, 56.16718,
    57.37427, 60.382, 62.78762, 62.45838, 64.11802, 70.75949, 69.12814,
    52.76382, 38.45281,
  78.4243, 81.85658, 83.97483, 85.42461, 87.27025, 86.56822, 75.7298,
    70.03649, 69.18489, 66.86583, 64.80667, 63.91088, 64.76899, 68.73979,
    70.13515, 64.75117, 65.10964, 66.42149, 65.08656, 61.58059, 60.54039,
    64.5013, 68.95971, 68.40401, 66.04662, 71.68504, 74.38441, 63.0755,
    42.1082, 39.30001,
  82.00832, 85.07242, 82.12497, 82.68536, 83.78798, 77.73997, 63.18715,
    67.9343, 68.9608, 71.96988, 75.42403, 79.10296, 78.79797, 77.40962,
    74.71799, 75.87201, 76.28583, 75.03362, 72.70808, 71.87638, 72.97254,
    71.94666, 69.62388, 65.45541, 69.31795, 77.16145, 70.36984, 48.79845,
    38.76358, 38.4239,
  81.44868, 82.14308, 83.27114, 83.80302, 87.74587, 82.16748, 75.07685,
    80.28942, 84.91495, 85.15815, 78.02613, 68.46612, 66.21519, 66.17801,
    65.82719, 66.29369, 66.70098, 66.34486, 66.32582, 68.21684, 72.09357,
    69.07973, 62.15178, 61.23817, 66.60809, 65.41364, 50.70258, 38.98844,
    39.3998, 38.3162,
  88.67709, 84.39303, 92.25141, 97.94167, 93.95073, 83.74864, 85.3884,
    79.48518, 73.8443, 71.4706, 65.89388, 62.4064, 64.13279, 64.10964,
    61.8297, 61.34555, 59.80092, 59.4273, 59.3828, 61.29776, 65.68793,
    64.98372, 61.05219, 66.63757, 67.52926, 54.03707, 39.90845, 41.62429,
    39.9588, 38.84364,
  108.8935, 111.7569, 114.0904, 113.8556, 111.745, 107.95, 92.50975,
    80.60324, 84.9984, 75.52155, 70.34147, 68.09557, 72.21431, 73.62038,
    67.90666, 58.88015, 59.68118, 59.10894, 58.84827, 61.21537, 64.61625,
    64.84885, 62.46184, 58.93181, 54.87349, 47.73539, 41.05106, 42.34328,
    41.20198, 39.72561,
  111.8822, 113.1872, 111.9817, 108.2382, 105.0226, 103.1403, 102.0111,
    100.8855, 94.83889, 93.74399, 97.10352, 93.69037, 91.29018, 89.58433,
    82.71727, 70.82877, 67.85715, 72.45373, 74.48853, 69.47659, 63.83387,
    59.6117, 54.15891, 47.46646, 43.33464, 42.43953, 41.07022, 40.42552,
    40.30978, 39.51314,
  106.4522, 101.613, 98.40681, 94.71893, 93.9247, 97.94183, 103.4071,
    101.4643, 95.04701, 94.17654, 89.90903, 84.64168, 83.79213, 85.45419,
    84.28203, 81.96664, 76.59364, 72.77829, 70.62847, 64.95617, 54.77931,
    51.36109, 45.51678, 42.31572, 42.04141, 41.60678, 40.63444, 39.69252,
    39.11611, 38.70774,
  91.65346, 91.89675, 91.92656, 90.65554, 89.36494, 90.32561, 91.1903,
    87.43753, 81.95001, 77.79596, 75.81285, 72.90461, 72.3963, 75.09864,
    72.12709, 69.84565, 68.12225, 62.50555, 58.30827, 52.9095, 46.60651,
    45.81693, 42.65118, 41.60516, 41.68761, 41.24493, 40.36795, 39.5858,
    38.98045, 38.60804,
  81.64801, 80.29944, 79.48276, 78.94254, 78.37712, 77.39419, 77.04056,
    77.12138, 74.90827, 71.30202, 67.19946, 69.82207, 73.72993, 70.40656,
    65.09779, 61.64096, 58.27525, 55.31174, 53.57515, 50.9007, 45.48002,
    45.36443, 42.89005, 41.66296, 41.47778, 41.28289, 40.1499, 39.09533,
    38.76105, 38.56021,
  71.07351, 71.33049, 70.44926, 70.93099, 71.20623, 71.82629, 72.3364,
    73.23843, 73.21453, 71.21822, 72.99743, 75.31786, 73.9799, 71.00173,
    65.3746, 60.30573, 55.74727, 54.39625, 54.67527, 51.39321, 45.28978,
    44.72116, 43.07769, 42.24129, 41.24513, 40.61152, 39.87953, 38.68194,
    38.50404, 38.39347,
  77.27892, 74.27705, 68.07117, 65.04773, 66.33055, 66.26521, 66.66,
    67.08522, 66.23965, 66.92722, 69.08556, 66.8976, 61.48815, 60.54344,
    58.92661, 59.72663, 63.76513, 67.46897, 66.1366, 60.31739, 51.53193,
    46.23193, 43.76536, 42.84865, 41.3512, 40.53601, 39.78607, 38.6799,
    38.45438, 38.39849,
  76.8046, 72.63808, 65.70479, 61.6253, 62.61286, 62.53438, 62.53212,
    62.51141, 63.32134, 66.02919, 66.14912, 61.80404, 61.03637, 59.79302,
    58.62003, 58.87608, 61.52929, 64.63652, 63.79581, 60.39862, 54.65308,
    48.94808, 45.24922, 43.99567, 42.70541, 41.07334, 40.03345, 38.90857,
    38.47332, 38.42176,
  74.36993, 70.78516, 63.67305, 60.29023, 61.11126, 61.28075, 61.42163,
    61.85876, 63.31232, 65.17661, 63.41027, 60.63774, 62.243, 61.0853,
    58.89758, 57.20979, 56.59005, 56.09128, 55.161, 53.26784, 51.89132,
    50.736, 47.87554, 45.88677, 43.95146, 41.62373, 39.92617, 38.99238,
    38.52518, 38.45169,
  72.40028, 69.73766, 63.70566, 61.22394, 61.80529, 61.14454, 61.69864,
    62.02874, 63.61196, 63.66374, 59.98165, 57.55388, 57.89375, 56.46847,
    54.53756, 53.09009, 51.68668, 50.84434, 50.73672, 50.61818, 50.43105,
    49.79858, 49.1725, 48.12397, 45.46744, 41.87608, 40.06145, 39.27206,
    38.61988, 38.4575,
  70.87802, 69.72614, 63.45962, 61.47374, 63.2186, 63.17165, 61.91033,
    59.88091, 59.46609, 57.64238, 54.02387, 53.49353, 53.35608, 52.62025,
    51.36258, 50.9695, 50.39004, 49.03024, 48.59116, 48.51218, 48.178,
    47.46988, 46.56585, 46.67659, 46.62722, 43.2444, 40.75543, 40.23015,
    39.24695, 38.50443,
  73.04411, 73.11263, 68.73444, 67.16544, 67.09106, 65.44673, 64.37794,
    62.95643, 63.29781, 60.48688, 57.48715, 58.72359, 59.39595, 58.92202,
    57.15967, 55.87759, 54.66399, 52.51875, 50.29321, 49.0365, 47.89622,
    47.25419, 46.22068, 45.82515, 46.55741, 46.08412, 43.57977, 41.29228,
    40.40383, 39.04796,
  75.37519, 72.87143, 67.61536, 65.25081, 64.51911, 63.01003, 63.29839,
    65.81166, 68.77253, 65.32103, 61.49483, 62.90036, 63.47976, 63.02904,
    61.34723, 60.18241, 58.12716, 55.93898, 53.4319, 51.53063, 50.41353,
    49.12933, 47.23008, 45.95131, 46.60542, 47.58084, 46.84768, 43.6499,
    41.77271, 40.05511,
  77.72594, 75.90579, 70.96722, 66.73677, 64.87857, 63.98409, 66.9558,
    71.22598, 71.29246, 66.74883, 65.67956, 66.22974, 66.52171, 65.02706,
    62.5363, 61.26326, 59.95856, 58.28749, 56.23902, 54.38917, 52.97832,
    51.25479, 48.22221, 46.59721, 46.87895, 47.05489, 47.18372, 44.73308,
    41.30916, 39.77264,
  79.20895, 76.49593, 71.6065, 68.20695, 66.67344, 65.34399, 68.52549,
    70.40942, 68.99438, 66.72772, 67.18855, 67.20343, 66.74319, 65.33485,
    63.05923, 61.4733, 60.31876, 59.16539, 57.44743, 56.10865, 55.98751,
    55.95023, 54.05686, 51.60929, 50.69915, 50.27271, 50.49105, 47.92252,
    41.87885, 38.85952,
  79.57668, 77.45943, 74.32192, 73.566, 73.85906, 72.83818, 72.66751,
    70.86175, 67.91293, 67.66061, 67.87319, 67.97282, 67.97316, 67.08345,
    65.49481, 63.76789, 62.49069, 61.64541, 60.86873, 60.53561, 59.48021,
    57.4572, 54.56573, 52.83671, 52.04429, 51.40132, 51.02353, 51.06968,
    47.3082, 40.5134,
  72.33414, 72.44391, 73.2068, 73.52705, 75.4245, 77.71637, 74.74677,
    68.04285, 65.48235, 65.44386, 64.59074, 64.23399, 64.60788, 64.92667,
    64.47487, 63.56959, 62.19145, 60.75822, 58.3008, 55.89859, 54.45397,
    52.60521, 50.38279, 49.0424, 48.759, 48.30781, 47.46623, 46.11779,
    44.78389, 41.43094,
  67.82854, 68.30653, 68.21351, 67.74619, 70.14716, 74.79088, 74.84919,
    67.64, 63.99712, 64.93871, 65.40247, 65.82972, 65.15437, 63.00687,
    60.27507, 57.67422, 54.1434, 51.16252, 49.93668, 48.30019, 46.90681,
    46.45002, 45.98523, 45.49662, 45.07731, 44.65779, 43.68934, 42.19144,
    40.4955, 38.77142,
  38.92716, 38.82604, 38.84991, 38.90849, 38.90985, 38.90943, 38.98627,
    39.16049, 39.40487, 39.79258, 40.49194, 40.39042, 39.2107, 39.44907,
    39.56857, 39.25265, 39.21344, 39.33004, 39.49416, 39.92128, 40.1413,
    39.59152, 39.67217, 40.6264, 41.91505, 42.36109, 43.54602, 45.05362,
    41.3487, 39.66495,
  39.48111, 39.47282, 39.25431, 39.52682, 39.43248, 39.3326, 39.55546,
    39.89133, 40.30638, 40.71163, 41.12522, 41.34507, 41.32061, 40.70458,
    40.23758, 40.34363, 39.71754, 39.86257, 40.14795, 40.29826, 40.02518,
    40.1649, 42.18848, 47.12259, 51.84648, 48.7364, 43.50161, 46.16965,
    41.89526, 40.16016,
  39.61443, 39.49342, 39.44061, 39.45897, 39.41655, 39.47119, 39.62975,
    39.8445, 40.05214, 40.23665, 40.4576, 40.7877, 41.05193, 41.30986,
    41.34672, 40.47954, 40.54123, 41.2317, 42.04163, 44.23908, 48.96497,
    55.77401, 60.46556, 61.50587, 60.05629, 54.40952, 50.02008, 45.69286,
    41.92055, 40.72076,
  39.5828, 39.58923, 39.9241, 40.34319, 40.74685, 41.27566, 41.36931,
    41.38871, 41.81665, 42.43124, 42.70436, 42.99735, 42.93246, 42.68121,
    43.99937, 44.98533, 44.87244, 45.78444, 49.8298, 56.02005, 64.55125,
    67.09598, 62.55814, 62.4531, 58.2303, 55.81955, 54.84226, 47.4773,
    41.04894, 39.6466,
  40.48542, 40.55205, 41.43612, 42.2637, 42.90887, 43.31053, 43.38098,
    43.19039, 43.23878, 42.61922, 41.26109, 40.70759, 40.9133, 42.37502,
    44.62051, 47.50784, 49.79024, 52.31524, 58.30999, 65.57757, 66.49547,
    57.61612, 53.27312, 55.085, 55.51855, 55.30265, 55.68595, 61.09939,
    59.81343, 46.60291,
  41.8115, 42.5593, 43.4659, 43.98325, 42.86216, 41.31088, 40.67624,
    40.08002, 40.53765, 42.58246, 46.82904, 56.54159, 66.80707, 67.24685,
    70.56413, 74.55386, 74.39233, 72.91788, 70.02803, 67.13579, 58.2906,
    48.82571, 51.79364, 54.52083, 58.22771, 60.68925, 63.8504, 75.08931,
    71.53455, 45.2303,
  42.27943, 42.5671, 43.05622, 43.69491, 44.14518, 46.98176, 55.07634,
    65.83591, 72.30688, 75.13222, 78.0941, 77.5538, 73.10938, 74.23848,
    75.32072, 75.30965, 74.55848, 68.46671, 61.28137, 57.52817, 52.52953,
    51.44738, 55.44802, 59.37305, 62.32237, 63.30351, 67.94283, 73.88116,
    61.22158, 38.93196,
  43.36611, 45.48391, 48.85938, 53.8275, 59.97413, 71.24694, 81.73538,
    77.34297, 73.77573, 74.20808, 71.34983, 67.02654, 63.46719, 62.57571,
    61.3005, 60.75956, 59.63734, 56.35215, 53.28004, 53.04271, 53.22497,
    55.07544, 58.38636, 61.35403, 61.77832, 63.48207, 69.35867, 68.05017,
    52.64282, 38.84991,
  52.33973, 57.43252, 62.56429, 68.27507, 75.51735, 80.04462, 72.6509,
    67.02808, 65.88369, 63.23723, 60.37677, 58.58212, 58.40634, 60.57034,
    61.04398, 56.71375, 57.03447, 58.87702, 59.11177, 57.28497, 56.957,
    60.33345, 64.33885, 64.69477, 63.687, 69.67526, 73.27328, 62.76712,
    42.20566, 39.47443,
  67.45267, 73.93947, 73.37386, 76.28488, 79.1977, 73.73135, 57.37471,
    59.42682, 58.63589, 59.821, 62.38533, 65.2378, 65.23886, 64.58662,
    62.78423, 64.13496, 65.94012, 66.32886, 65.75558, 65.42831, 66.6901,
    66.69672, 65.74014, 63.14773, 67.23209, 75.62155, 70.47908, 49.18542,
    38.98298, 38.99869,
  74.75993, 77.33409, 76.37621, 74.10822, 75.17331, 66.96785, 58.77557,
    64.16012, 68.52467, 70.72273, 66.62115, 59.66071, 58.24257, 58.49461,
    58.72495, 60.47155, 61.74907, 62.30099, 63.30556, 65.4896, 69.18984,
    67.40865, 62.25973, 62.48131, 69.1414, 68.397, 52.27985, 39.27906,
    39.60669, 38.83844,
  76.84301, 68.91795, 71.60987, 74.8896, 72.71689, 66.56503, 71.88708,
    68.93658, 64.46758, 64.20118, 58.86497, 55.27477, 57.36817, 57.82446,
    56.59765, 57.9234, 57.83484, 58.47197, 59.09366, 60.89267, 64.6387,
    64.20705, 61.15851, 66.31471, 68.36771, 55.84471, 39.90244, 41.14735,
    40.13992, 39.20697,
  87.49644, 88.76972, 91.84705, 93.44579, 93.60146, 91.71732, 80.48448,
    67.59834, 72.66391, 65.2613, 60.56973, 60.33432, 64.84158, 66.62389,
    62.92805, 55.45111, 56.66678, 56.99506, 57.31334, 59.48674, 63.25491,
    64.71538, 63.31335, 59.60172, 54.71784, 47.339, 40.39365, 42.14489,
    41.06599, 39.979,
  93.0319, 96.20294, 97.00504, 94.45496, 91.34563, 87.88933, 84.9656,
    84.25584, 79.62869, 79.17001, 83.56222, 82.20575, 80.70662, 80.27261,
    73.87126, 63.06601, 61.94547, 67.50471, 71.36911, 68.27728, 64.7905,
    61.10745, 54.93235, 48.12304, 43.38171, 42.15105, 41.07809, 40.77048,
    40.48962, 39.87331,
  94.84787, 94.25525, 90.96204, 87.25237, 83.55087, 84.06999, 85.89481,
    85.97764, 84.43895, 84.19789, 82.04353, 76.44827, 75.59923, 77.58704,
    77.62151, 76.67582, 73.19499, 72.167, 71.08987, 66.01105, 56.57296,
    52.28959, 45.54851, 41.98564, 41.80731, 41.52417, 40.76663, 39.97757,
    39.53127, 39.17731,
  90.57162, 87.47685, 84.17101, 81.73579, 81.41878, 83.90236, 85.23273,
    81.55679, 76.71629, 72.12672, 69.56888, 67.52499, 68.25835, 72.27805,
    71.03941, 69.3791, 68.02864, 63.18943, 58.71499, 53.20355, 47.10233,
    45.25568, 42.0085, 41.30859, 41.70766, 41.36074, 40.50621, 39.80898,
    39.31155, 39.04062,
  81.00591, 78.46639, 77.8445, 77.33986, 76.28015, 74.09956, 72.34576,
    71.51167, 68.71951, 65.60558, 63.20151, 66.10759, 70.40729, 68.54065,
    63.6137, 60.36154, 57.26633, 54.0878, 51.73886, 48.93298, 44.25481,
    43.87486, 41.92164, 41.21301, 41.39795, 41.39406, 40.38848, 39.49308,
    39.18714, 39.03525,
  72.76035, 72.47888, 70.83924, 69.52433, 67.57832, 66.37479, 66.12009,
    66.79716, 66.76892, 65.69948, 67.68568, 70.53025, 70.03235, 66.84369,
    61.05436, 56.28688, 52.1535, 50.52021, 50.35125, 47.81834, 43.4115,
    43.45512, 42.17517, 41.61062, 41.19843, 40.85442, 40.19189, 39.19995,
    39.01721, 38.91066,
  77.12845, 73.07391, 66.23029, 62.15128, 62.51473, 62.35946, 62.97866,
    63.66531, 63.25219, 63.87872, 65.45163, 63.22786, 57.63612, 55.30989,
    52.37335, 51.85671, 54.69269, 58.34592, 58.75654, 55.34135, 49.13464,
    45.22535, 42.96801, 42.35116, 41.29655, 40.81386, 40.22178, 39.2,
    38.94754, 38.88787,
  75.78893, 70.01524, 62.9528, 58.8064, 59.72134, 59.53105, 59.4128,
    58.95383, 58.75652, 59.82382, 58.77441, 54.02721, 52.21938, 50.89446,
    50.10645, 51.34628, 55.30029, 59.83002, 60.36163, 57.69159, 52.66083,
    47.52186, 44.29297, 43.55727, 42.4396, 41.25254, 40.41719, 39.39671,
    38.94867, 38.91423,
  71.93127, 67.15036, 60.12792, 56.23471, 56.27555, 55.51193, 54.74144,
    54.13526, 54.25755, 54.92514, 53.17264, 50.85234, 53.10191, 53.62782,
    53.5645, 54.1013, 55.4062, 55.96955, 54.8012, 52.03491, 49.85115,
    48.50421, 46.59574, 45.28108, 43.553, 41.71305, 40.36423, 39.45901,
    38.97227, 38.92736,
  68.57845, 64.50895, 57.65559, 53.85452, 53.35117, 52.04109, 52.01437,
    52.17344, 53.60366, 54.44914, 52.71027, 52.07857, 53.99057, 54.23697,
    53.58929, 52.86859, 51.72213, 50.58211, 49.60753, 48.69672, 48.26772,
    48.08231, 48.07099, 47.03619, 44.76458, 41.86367, 40.36262, 39.62714,
    39.06879, 38.94921,
  65.55122, 62.70525, 55.30079, 52.30852, 53.34629, 53.40246, 53.1595,
    52.56288, 53.26406, 52.94727, 51.12242, 51.17858, 51.45536, 50.99223,
    49.82934, 49.19201, 48.52488, 47.51303, 47.18092, 47.16343, 47.13174,
    46.93708, 46.31741, 45.79013, 45.32916, 42.55048, 40.59484, 40.24454,
    39.54203, 39.00154,
  65.78065, 64.34814, 59.15789, 57.28611, 57.62875, 56.71114, 56.52135,
    56.03733, 57.03618, 55.18763, 52.82238, 53.56224, 54.3047, 54.04617,
    52.71704, 51.98814, 51.39352, 50.21153, 48.6729, 47.73293, 47.12012,
    46.72629, 45.63974, 44.90455, 45.2929, 44.70942, 42.77867, 41.09823,
    40.44146, 39.46176,
  68.09804, 65.33559, 59.67417, 57.03534, 56.53488, 55.26967, 55.57823,
    57.56385, 60.17384, 57.59264, 54.58312, 56.06651, 57.38197, 57.56147,
    56.28568, 55.79233, 54.90648, 53.45304, 51.41255, 49.82486, 49.12103,
    48.14265, 46.23569, 44.97037, 45.52384, 46.18744, 45.56188, 43.03833,
    41.59041, 40.29516,
  68.4526, 65.97813, 60.87414, 56.96357, 55.72994, 54.92141, 57.17234,
    60.7057, 61.35517, 57.73751, 57.1431, 58.50542, 59.81945, 59.38964,
    57.66747, 57.15002, 56.68571, 55.61392, 53.85789, 52.33337, 51.25397,
    49.69074, 47.0142, 45.59528, 46.02307, 46.17688, 46.24333, 44.35063,
    41.50349, 40.18311,
  68.36096, 65.74056, 60.79801, 57.18691, 56.32109, 55.44065, 57.99675,
    60.07393, 59.62634, 57.89433, 58.73124, 59.79665, 60.43973, 59.7161,
    58.19757, 57.53168, 56.92395, 56.12038, 54.85649, 53.75899, 53.15793,
    52.60997, 50.93581, 49.13541, 48.63372, 48.43052, 48.62557, 46.75652,
    41.79149, 39.35973,
  68.2016, 65.58502, 61.95842, 60.68578, 61.3286, 60.85232, 61.32256,
    60.60272, 58.83187, 58.94772, 59.62378, 60.44965, 61.20479, 61.07075,
    60.25763, 59.25207, 58.4906, 58.20134, 58.10727, 58.17617, 56.78689,
    54.66982, 52.16563, 50.71586, 50.17902, 49.64881, 49.22728, 48.8149,
    45.49325, 40.43567,
  62.05023, 61.6747, 61.77069, 61.87593, 63.40888, 65.12444, 62.98488,
    58.60913, 57.06052, 57.40488, 57.10968, 57.40917, 58.50986, 59.56898,
    59.923, 59.69441, 59.16806, 58.53944, 57.04249, 55.38476, 53.81858,
    52.00666, 50.15253, 48.96436, 48.69395, 48.11797, 47.15068, 45.7171,
    44.12157, 41.28881,
  58.54086, 58.93781, 59.11092, 58.69177, 60.56634, 64.13422, 64.2146,
    58.74771, 56.29932, 57.24485, 57.94191, 59.04195, 59.49948, 58.76049,
    57.26846, 55.75558, 53.54021, 51.54245, 50.47286, 49.08741, 47.78862,
    47.20676, 46.76478, 46.19931, 45.69727, 45.13717, 43.95422, 42.36776,
    40.9747, 39.39047,
  5.344968, 4.568901, 4.894967, 5.01931, 5.11331, 5.23462, 5.445849,
    5.724692, 6.169326, 7.00659, 8.610914, 10.53384, 11.9932, 15.07352,
    18.67568, 22.74639, 27.45251, 33.02921, 38.88509, 44.18027, 48.92573,
    52.05158, 54.05939, 55.5748, 55.55822, 53.21615, 51.53066, 54.02779,
    48.38901, 46.26052,
  4.473154, 3.937462, 4.132336, 4.638041, 4.912834, 5.12639, 5.485184,
    5.723316, 6.018306, 6.584429, 7.848266, 10.06077, 12.91366, 15.46845,
    18.72115, 23.52768, 29.22425, 35.52307, 40.31106, 45.51828, 50.12085,
    54.10408, 56.96436, 58.83607, 59.56656, 58.87878, 51.2091, 52.48583,
    48.62919, 46.87333,
  6.996668, 6.927335, 7.786894, 8.352596, 9.068319, 9.939159, 10.69449,
    11.38055, 11.86708, 12.17469, 12.5795, 13.51004, 15.15196, 17.51687,
    20.33951, 23.09822, 28.06917, 35.18849, 41.39703, 46.88477, 52.10051,
    56.32964, 59.1011, 60.37946, 60.41053, 59.82344, 59.32135, 53.72871,
    47.75505, 46.83454,
  9.69546, 10.17574, 11.48123, 12.41525, 13.00332, 13.8248, 14.56759,
    15.59821, 16.20556, 16.76764, 17.77384, 19.08798, 20.78275, 22.91476,
    25.39716, 28.14116, 30.81754, 34.69312, 41.40527, 46.9643, 52.38985,
    56.6554, 58.89573, 60.53973, 60.68808, 60.6692, 60.63478, 59.57341,
    55.32137, 47.41097,
  12.169, 12.97309, 14.69316, 15.80924, 15.89113, 15.89127, 15.96787,
    16.03396, 16.35167, 17.12443, 18.38976, 20.1887, 22.20827, 24.55696,
    27.2862, 30.41531, 33.92596, 37.85435, 42.51269, 47.99688, 52.74728,
    56.00218, 58.61593, 60.09576, 60.51357, 60.5176, 60.26071, 61.04018,
    60.62294, 56.96619,
  11.74183, 13.18493, 15.43694, 16.35643, 16.43814, 16.44089, 16.67612,
    16.82501, 16.84103, 17.20969, 18.27813, 20.10157, 22.69642, 25.1774,
    28.1435, 31.61688, 35.69545, 39.88688, 44.29748, 49.26328, 53.4212,
    54.1499, 58.95948, 60.12641, 60.36262, 60.03537, 59.51976, 60.11861,
    60.08999, 50.93036,
  11.95883, 12.81447, 14.76573, 16.3046, 16.59019, 16.88623, 17.3295,
    17.77576, 18.03913, 18.34249, 19.09205, 20.08182, 17.27108, 20.98893,
    25.15116, 30.56106, 34.60569, 39.25673, 43.82619, 49.15263, 53.59492,
    57.00447, 59.31207, 60.49114, 60.49463, 59.82823, 59.68801, 59.78937,
    59.06894, 44.94147,
  16.86097, 15.9423, 16.38417, 16.47786, 16.62461, 17.0848, 17.47401,
    16.04956, 11.72751, 15.05721, 16.45283, 17.33584, 19.51777, 22.84499,
    26.61745, 30.53256, 34.85207, 39.56291, 44.38832, 49.37888, 53.95963,
    57.40287, 59.65134, 60.58294, 60.33551, 60.10609, 60.24572, 59.78227,
    58.09091, 45.18536,
  19.68553, 17.97933, 17.76973, 17.50982, 17.33262, 17.25513, 16.25924,
    13.40906, 13.74311, 14.30905, 16.38797, 18.95267, 22.12119, 25.06027,
    28.26047, 30.91133, 34.93965, 40.28591, 45.68948, 50.45803, 54.74064,
    58.14426, 60.03691, 60.46511, 60.09777, 60.39444, 60.33181, 59.27612,
    45.4483, 45.76715,
  24.74097, 22.66999, 21.185, 20.09385, 19.60124, 18.64371, 16.72886,
    17.01487, 16.95679, 17.52886, 18.20107, 20.91747, 23.28468, 25.05232,
    27.19545, 31.1557, 35.21279, 39.96658, 45.23912, 50.73152, 55.66703,
    58.56933, 59.50711, 59.3478, 59.68299, 60.03317, 59.53802, 51.69517,
    45.13189, 44.8559,
  29.78169, 27.12129, 26.98938, 24.49261, 23.26341, 21.40286, 19.78248,
    18.81308, 18.52467, 19.22495, 19.93732, 21.34001, 22.96773, 23.78768,
    25.67034, 29.31817, 33.48248, 38.64461, 44.3727, 49.60079, 55.14837,
    58.29929, 59.06981, 59.2873, 59.69361, 59.31235, 53.42343, 45.4461,
    46.01691, 44.93137,
  30.46218, 28.20758, 30.80297, 30.90267, 29.50941, 25.77713, 22.47615,
    19.58348, 18.4712, 18.95103, 20.05813, 21.66626, 24.21666, 26.2993,
    28.62902, 32.04544, 35.37202, 38.78034, 42.65821, 48.26133, 54.17072,
    57.90978, 58.82236, 59.59861, 59.86572, 58.85746, 45.75185, 49.58354,
    46.52429, 45.59132,
  20.52727, 22.00998, 24.3293, 27.23511, 29.44226, 28.99384, 22.6795,
    17.34949, 20.8946, 19.71345, 21.1658, 22.22342, 24.30351, 26.62341,
    29.16909, 31.55939, 35.59111, 40.02374, 44.89377, 49.84549, 54.29791,
    57.28689, 58.57565, 55.27285, 55.00896, 53.91053, 46.37601, 47.89012,
    47.42752, 46.31789,
  16.60934, 15.51172, 15.64401, 15.89527, 16.45874, 17.24707, 18.20529,
    19.46428, 18.36714, 19.51771, 21.3417, 23.31484, 25.05067, 26.8831,
    29.585, 32.21987, 35.16864, 40.38102, 45.65176, 50.34797, 53.90494,
    56.55973, 53.50723, 48.90795, 46.05864, 46.30235, 45.83724, 45.43634,
    45.64238, 45.69784,
  17.46264, 11.349, 14.63332, 15.15452, 17.09539, 17.38108, 17.72972,
    17.89689, 18.29362, 19.4948, 21.10799, 23.02652, 25.12871, 27.39876,
    29.3122, 31.94525, 35.77122, 39.07408, 44.5901, 49.78067, 48.72221,
    51.56386, 49.38569, 47.24407, 47.54784, 46.81278, 46.15472, 45.63446,
    45.16864, 45.05644,
  9.50313, 10.82817, 12.60074, 14.63771, 16.51638, 17.63976, 18.27158,
    18.60096, 19.09544, 20.59247, 22.73628, 24.50004, 26.36316, 27.97548,
    29.88613, 32.52142, 35.39931, 38.94131, 39.9761, 43.86824, 44.54199,
    47.9062, 47.71979, 47.41338, 47.30433, 46.74746, 46.12645, 45.69608,
    45.22723, 45.07535,
  6.994177, 5.594076, 7.11941, 8.6309, 10.38831, 12.67411, 15.17211,
    17.77596, 18.94523, 20.6661, 22.60452, 25.31257, 28.43326, 30.15339,
    32.10018, 34.22975, 36.7611, 40.12148, 42.6257, 45.41268, 44.9598,
    47.97305, 47.93997, 47.41803, 47.32969, 46.93052, 45.98446, 45.21099,
    44.9553, 44.97013,
  10.37948, 7.319107, 6.24566, 6.494779, 7.66285, 8.78141, 10.16319, 11.6725,
    14.00285, 16.5684, 21.09858, 24.18178, 27.02182, 30.84476, 33.99105,
    36.42345, 39.07642, 43.22414, 48.24676, 51.40848, 48.02606, 48.42543,
    48.10624, 47.75338, 47.09894, 46.65551, 46.05827, 45.07779, 44.83175,
    44.87019,
  24.05384, 16.58257, 9.268264, 4.047017, 6.02152, 6.162177, 7.120747,
    8.109665, 9.20216, 11.26445, 14.55543, 17.24329, 19.17834, 24.70376,
    31.14541, 35.99022, 40.3469, 45.82856, 51.60265, 55.8364, 56.86818,
    52.43793, 49.69869, 49.32241, 47.98714, 47.08409, 46.32926, 45.26554,
    44.81851, 44.90223,
  23.38904, 16.86579, 9.555536, 4.550473, 5.965967, 6.15703, 7.038429,
    8.084213, 9.792987, 12.54883, 14.74246, 14.92649, 17.70185, 19.94982,
    23.21259, 27.49429, 33.53289, 41.07223, 48.19691, 53.50758, 56.15212,
    55.15205, 52.03895, 50.87725, 49.38115, 47.75006, 46.64643, 45.46137,
    44.7952, 44.91372,
  25.47109, 18.95956, 11.67319, 6.763876, 7.659576, 7.51753, 8.10731,
    8.915428, 10.46953, 12.3643, 13.29284, 14.13907, 18.0073, 20.724,
    23.32979, 26.97004, 31.82289, 37.82283, 43.90204, 48.65602, 52.38482,
    55.01702, 54.5105, 52.68476, 50.63599, 48.39222, 46.79059, 45.48588,
    44.78798, 44.91847,
  27.85159, 22.20195, 15.27605, 11.33002, 12.72774, 12.10488, 12.51816,
    12.76698, 14.16759, 15.35457, 15.19387, 16.38309, 19.46178, 22.31814,
    25.07013, 28.80017, 33.19532, 38.19473, 43.40266, 47.59463, 50.91962,
    53.02101, 54.43337, 54.42223, 52.56404, 49.39802, 47.26677, 45.97102,
    44.91008, 44.89478,
  28.71246, 24.63024, 18.35777, 15.13085, 17.78386, 18.64853, 19.20117,
    18.95193, 19.53038, 20.0501, 20.53045, 23.2007, 25.97627, 28.57359,
    30.87176, 34.24067, 38.16333, 41.80861, 45.66629, 48.87393, 51.35935,
    52.88366, 53.38068, 53.6116, 53.88554, 51.2498, 48.33268, 46.79643,
    45.70842, 45.0421,
  29.07965, 25.163, 20.04433, 17.91406, 19.96288, 20.61637, 22.48552,
    24.09626, 25.84014, 25.65725, 26.38939, 30.7645, 35.01667, 38.13902,
    39.89159, 42.53418, 45.66439, 48.63464, 51.24901, 53.70626, 55.41501,
    55.69044, 54.97785, 54.24604, 54.52157, 54.09087, 51.42588, 48.08139,
    46.78534, 45.77246,
  28.91076, 23.9678, 18.25936, 15.13514, 17.18923, 18.32051, 20.0205,
    22.69837, 25.29739, 25.64119, 25.81313, 30.00578, 34.57427, 38.14811,
    40.11153, 43.24855, 46.11945, 49.49458, 52.92417, 55.93211, 57.89366,
    57.95106, 56.08006, 54.36932, 54.33029, 54.01987, 53.0108, 49.72173,
    47.38947, 46.47361,
  30.34805, 26.48742, 21.16406, 17.18199, 17.96326, 18.66637, 21.35905,
    24.36271, 25.08318, 25.5977, 27.96213, 31.5002, 35.72795, 38.41347,
    39.82773, 42.51712, 45.56297, 48.58062, 52.58835, 56.51059, 59.23257,
    60.12124, 58.2867, 56.26509, 55.81828, 54.74769, 53.97264, 50.99586,
    46.9351, 45.98681,
  37.1487, 33.66509, 28.15935, 24.34163, 24.86136, 24.6895, 26.80361,
    28.19288, 28.41466, 29.55949, 32.75695, 36.24215, 39.82336, 42.07578,
    43.04637, 44.96092, 46.77079, 49.02797, 52.41007, 55.78949, 58.39772,
    60.10633, 59.53354, 58.08627, 57.59698, 56.87352, 56.47733, 54.0787,
    48.59948, 45.55558,
  47.50616, 45.82521, 41.84077, 40.01161, 40.95164, 40.43368, 39.75937,
    38.95101, 37.87506, 38.74245, 40.18853, 42.66151, 45.64693, 47.43556,
    48.00289, 48.82368, 49.21913, 50.19134, 52.45634, 55.12358, 56.10187,
    56.06832, 54.91761, 54.042, 54.32106, 54.10788, 53.66531, 53.56593,
    51.65892, 46.94075,
  46.89553, 47.56529, 49.18171, 51.1005, 52.50815, 53.79836, 51.81254,
    47.59565, 46.39336, 46.90162, 46.71026, 46.87785, 47.29529, 47.95687,
    48.22309, 48.38989, 48.2223, 48.24028, 48.5928, 48.9675, 49.83643,
    50.78908, 50.76181, 50.08707, 50.25377, 50.23316, 49.62201, 48.30102,
    47.88633, 47.09905,
  49.11254, 49.82054, 50.05947, 49.95752, 51.21417, 53.67664, 54.1071,
    50.81571, 48.63205, 49.43465, 49.95739, 50.54745, 50.70245, 50.19994,
    49.64088, 49.03233, 47.81773, 46.52275, 46.38804, 46.51302, 46.292,
    46.94011, 47.75559, 48.14482, 47.99516, 48.23782, 47.97652, 46.83534,
    45.88715, 45.10409,
  26.08447, 28.23257, 30.60328, 33.26056, 35.78152, 38.15662, 40.69003,
    43.35561, 46.15936, 49.06824, 51.97423, 54.57019, 56.57346, 58.19577,
    59.41656, 60.25334, 60.82288, 61.39027, 61.98945, 62.74599, 63.56174,
    64.38659, 65.39163, 66.35047, 66.94897, 65.99295, 57.44642, 60.36081,
    56.08817, 53.62806,
  26.67416, 28.28281, 30.6533, 33.04599, 35.57352, 38.29435, 41.05597,
    43.88557, 46.77311, 49.66769, 52.5462, 55.32285, 57.64525, 59.1409,
    59.98729, 60.59201, 60.95404, 61.42594, 62.12755, 63.10083, 64.25229,
    65.48666, 66.74929, 68.01784, 68.88403, 68.24636, 64.74109, 58.41999,
    55.37389, 53.89179,
  27.37751, 28.86506, 31.28267, 33.57732, 35.99266, 38.76646, 41.61104,
    44.66693, 47.77357, 50.64095, 53.3888, 55.97734, 58.27986, 59.98254,
    60.96476, 61.29668, 61.40751, 61.67338, 62.23167, 63.04976, 64.46198,
    66.10983, 67.45181, 68.64273, 69.21262, 69.42078, 68.86756, 67.05571,
    55.61687, 53.49604,
  27.83713, 29.48877, 31.95959, 34.29068, 36.60783, 39.04433, 41.68678,
    44.72795, 47.92612, 51.12622, 54.05924, 56.59795, 58.8837, 60.50996,
    61.62852, 62.24345, 62.17805, 62.07947, 62.5934, 63.39583, 64.56305,
    65.64413, 66.24367, 67.85015, 68.61909, 69.46455, 69.9555, 69.13834,
    67.2228, 56.00567,
  28.37332, 30.0475, 32.71306, 35.17688, 37.55722, 39.78557, 42.08175,
    44.94934, 47.80379, 50.97933, 54.04348, 56.86075, 59.50025, 61.27546,
    62.40881, 63.08776, 63.1935, 62.9824, 63.16356, 63.89941, 64.44242,
    64.60257, 65.89513, 67.3205, 68.35126, 68.88409, 69.1076, 70.21188,
    69.7749, 66.84293,
  29.16364, 30.53122, 33.07055, 35.68941, 38.25926, 40.63243, 42.86474,
    45.94714, 48.50941, 50.9145, 53.68781, 56.4883, 59.43513, 61.34826,
    62.70821, 63.58726, 63.80716, 63.81078, 63.62427, 63.93369, 64.14138,
    64.39002, 66.16203, 67.5695, 68.35079, 68.56465, 68.39358, 69.05696,
    69.05773, 58.34705,
  32.07713, 32.26063, 34.20629, 36.15979, 38.61078, 41.10748, 43.54321,
    46.55193, 49.41564, 51.77119, 54.19569, 56.00256, 57.23676, 59.28171,
    60.76116, 61.85621, 62.53265, 62.68467, 62.48848, 62.92636, 63.49374,
    64.50163, 66.05785, 67.65466, 68.47418, 68.51756, 68.61062, 68.63918,
    67.80045, 52.13899,
  37.4899, 36.51003, 37.16417, 38.0654, 39.76299, 42.20542, 44.63589,
    45.70399, 47.57479, 50.17992, 52.54842, 54.70119, 56.89222, 58.99797,
    60.57463, 61.5682, 62.555, 63.21759, 63.23482, 63.29702, 63.74194,
    64.62427, 65.96236, 67.31752, 68.05421, 68.67954, 69.04098, 68.44237,
    66.74866, 52.46265,
  43.67494, 43.43246, 42.57025, 42.27318, 42.66928, 44.01424, 44.43685,
    46.39646, 48.86797, 51.0974, 53.21172, 55.11436, 56.85453, 58.81549,
    60.61741, 61.24732, 62.15081, 63.44281, 64.37473, 64.43488, 64.62062,
    65.13638, 65.9531, 66.79601, 67.54636, 68.57367, 68.95356, 67.87249,
    52.3802, 53.06855,
  46.47867, 49.11982, 49.43968, 48.4635, 47.49982, 46.8539, 46.12275,
    47.86884, 49.83749, 52.18184, 54.01325, 55.86238, 57.32162, 58.50872,
    59.49792, 60.66626, 61.58821, 62.56034, 63.52373, 64.21501, 65.10411,
    65.30785, 65.66547, 66.222, 67.37446, 68.03631, 67.76155, 59.64304,
    52.84785, 52.21922,
  44.35191, 47.48892, 52.21802, 53.71915, 53.41005, 51.2824, 49.93836,
    50.26505, 51.13705, 53.61298, 55.10971, 56.19, 57.37821, 58.44056,
    59.40812, 60.24611, 61.03411, 61.37856, 61.0553, 62.22661, 64.42556,
    64.8161, 65.06583, 66.39045, 67.9521, 67.67691, 63.25113, 54.06425,
    53.76647, 52.51733,
  40.25529, 40.25321, 47.86576, 53.52122, 58.12842, 56.58596, 53.02543,
    50.82865, 52.31041, 53.57262, 55.62908, 56.91109, 58.7216, 59.63081,
    59.98698, 60.37096, 61.17614, 61.91847, 62.60638, 62.66096, 64.03211,
    64.6018, 64.63567, 66.06533, 67.65096, 67.23655, 52.55469, 58.39442,
    54.75242, 53.30793,
  33.87395, 36.39215, 39.19178, 44.89639, 51.44666, 56.29979, 53.66954,
    49.32212, 54.97097, 55.22002, 57.33142, 58.62142, 60.20379, 61.36783,
    61.6824, 60.53953, 61.29917, 62.33497, 63.13964, 63.39632, 64.05943,
    64.56754, 64.80573, 60.61203, 60.13314, 62.47194, 53.17592, 54.63489,
    55.05573, 54.05596,
  32.4219, 34.00334, 35.61777, 37.77176, 39.85095, 43.39943, 47.73619,
    52.30673, 52.91758, 55.58945, 58.17958, 60.37169, 61.59391, 62.52945,
    62.7789, 61.98304, 61.31821, 62.13883, 63.34275, 63.38827, 63.34061,
    63.92772, 60.74798, 55.55451, 52.3628, 53.11412, 53.36205, 52.4712,
    52.6548, 53.02243,
  30.56323, 26.76923, 34.5827, 37.77733, 40.73048, 43.7373, 46.3162,
    49.16793, 52.69521, 55.58175, 57.86706, 59.76113, 61.56944, 63.05772,
    63.41493, 63.64368, 62.78418, 61.78254, 61.7061, 62.13948, 57.29779,
    58.21582, 55.6885, 53.31483, 54.54808, 54.07916, 53.5636, 53.01359,
    52.49227, 52.40033,
  23.37295, 25.57245, 28.23762, 31.85664, 35.93863, 40.96491, 44.78475,
    47.74365, 50.93095, 54.45755, 57.35531, 59.59327, 61.53817, 63.32628,
    64.12127, 64.31512, 64.30617, 63.23355, 60.64065, 57.24373, 54.1847,
    55.12768, 54.15372, 53.7097, 54.05477, 53.91521, 53.27431, 52.82545,
    52.54098, 52.44601,
  27.5674, 25.72603, 28.52318, 31.01936, 33.75654, 37.10543, 40.91935,
    44.91487, 49.71602, 52.80532, 55.61888, 58.63243, 61.34761, 62.91316,
    64.09897, 65.06895, 65.65384, 65.65365, 64.89767, 63.20975, 56.00117,
    55.44926, 54.66233, 54.14665, 54.45751, 54.36373, 53.33583, 52.49274,
    52.29434, 52.30191,
  39.0036, 33.33324, 31.49131, 32.45748, 35.94613, 38.54589, 41.68148,
    44.87923, 48.03294, 50.79543, 55.12564, 58.20716, 60.01668, 61.67668,
    62.86464, 64.10795, 65.49632, 66.85212, 67.62514, 66.99253, 62.77258,
    57.28756, 55.31857, 55.32602, 54.72408, 54.6325, 53.80306, 52.4899,
    52.25058, 52.21264,
  51.00034, 46.34425, 39.37955, 33.43637, 37.96964, 40.04875, 43.2932,
    46.31391, 49.39009, 52.54809, 55.9158, 57.38716, 56.55699, 56.7472,
    57.82848, 59.96626, 63.91607, 65.84889, 67.44118, 68.44422, 68.01075,
    63.33016, 57.79852, 57.66916, 56.2458, 55.44821, 54.46774, 52.79016,
    52.21136, 52.26524,
  50.18818, 47.09071, 41.89988, 37.16615, 40.96189, 43.05322, 46.347,
    49.40698, 52.73422, 56.08046, 58.80735, 59.75598, 61.8409, 60.36553,
    59.14391, 58.4353, 59.02058, 61.1132, 62.99751, 64.88081, 66.76254,
    65.76106, 61.41659, 59.84324, 58.29811, 56.43708, 54.77294, 53.13355,
    52.14523, 52.28872,
  51.62, 48.35392, 44.61454, 40.91822, 44.7831, 46.70541, 49.89845, 53.28874,
    56.8983, 59.78248, 60.924, 61.05316, 63.36246, 64.02835, 62.88029,
    62.57281, 62.29573, 62.78547, 62.69479, 61.94817, 62.34356, 63.85987,
    63.98096, 62.33291, 60.62288, 57.61492, 55.32069, 53.20636, 52.18362,
    52.28513,
  54.47862, 51.22427, 47.30598, 45.05279, 49.24935, 51.35517, 54.31393,
    57.22282, 60.52707, 63.62956, 65.86915, 67.33583, 68.48521, 68.74687,
    67.82804, 66.77317, 65.88541, 65.30175, 64.7187, 63.45102, 62.58281,
    62.09485, 63.2047, 63.36353, 62.55676, 59.26612, 56.05999, 54.10484,
    52.55434, 52.24346,
  59.61522, 56.83092, 52.58316, 50.19779, 53.52742, 55.37726, 58.0789,
    60.73508, 63.5696, 66.45947, 69.25091, 71.95326, 73.79819, 74.30599,
    73.66961, 72.7914, 71.81382, 70.79925, 69.05877, 67.15215, 65.6914,
    64.17902, 63.24012, 62.9698, 63.61866, 61.12292, 57.32377, 55.34512,
    53.7229, 52.58839,
  67.16045, 63.22049, 58.73106, 56.25555, 58.30612, 59.3007, 61.55947,
    64.26795, 67.14077, 69.25195, 71.51946, 75.08323, 78.44265, 79.96538,
    79.33855, 78.63882, 77.19646, 75.51198, 73.98699, 72.80773, 71.34778,
    69.02229, 66.2754, 64.64638, 64.66885, 63.78073, 60.66728, 56.71794,
    55.03672, 53.61893,
  73.38156, 68.7878, 63.27161, 57.98813, 59.797, 60.46938, 62.97421,
    65.64735, 68.33252, 69.64851, 71.10345, 73.81532, 77.30953, 78.99512,
    78.46727, 78.4977, 77.69443, 76.2681, 74.42297, 73.42367, 72.84579,
    71.07649, 67.53341, 65.48154, 65.36488, 64.23015, 62.3354, 58.10507,
    55.14175, 54.20037,
  77.00866, 71.96567, 66.84312, 61.41669, 61.69406, 61.2156, 63.59863,
    66.50034, 68.22415, 68.49927, 70.59097, 73.66347, 76.69064, 78.00398,
    77.26553, 77.06903, 76.70095, 75.05689, 73.0724, 72.32918, 71.91515,
    70.99919, 68.06238, 65.92631, 65.95424, 65.02042, 63.82365, 60.02682,
    55.02182, 53.57627,
  77.68056, 74.06112, 69.12364, 63.95553, 64.13784, 62.36834, 63.25397,
    64.54333, 64.86034, 64.94321, 67.01266, 70.50929, 74.20403, 75.61813,
    74.12403, 73.84336, 72.99944, 72.12154, 71.2435, 70.57635, 70.04225,
    69.31759, 67.24452, 65.21597, 65.12229, 64.72367, 64.53677, 62.68259,
    57.33884, 53.40384,
  73.97756, 71.89949, 68.09887, 65.498, 66.66888, 65.62193, 64.01972,
    63.06165, 62.12853, 62.10062, 62.55769, 64.4858, 67.59922, 68.87082,
    67.91381, 67.51983, 66.43217, 65.57832, 65.66995, 66.39058, 66.4097,
    65.57829, 63.10915, 61.54182, 61.84204, 61.42848, 60.5712, 60.1344,
    58.88923, 54.71259,
  59.1904, 60.14452, 61.54344, 63.11824, 64.25659, 65.8737, 63.75342,
    59.86836, 58.41565, 59.00636, 58.71577, 58.73932, 58.77982, 59.32082,
    58.81165, 58.60717, 57.89336, 57.18512, 56.73437, 56.59074, 57.077,
    58.44669, 58.80605, 58.12814, 58.42238, 58.52584, 57.67681, 55.54522,
    54.63322, 54.30777,
  56.24256, 56.93858, 57.40102, 57.10124, 57.87037, 59.5878, 60.44129,
    57.62621, 55.6622, 56.11744, 56.43954, 56.96447, 57.09164, 56.61209,
    56.14377, 55.65327, 54.75367, 53.66341, 53.47266, 53.45235, 53.13418,
    53.72116, 54.73305, 55.44543, 55.42019, 55.58578, 55.44524, 54.25098,
    53.09123, 52.41553,
  57.75857, 59.31488, 60.48109, 61.54353, 62.4548, 63.24373, 63.89169,
    64.40114, 64.82361, 65.29742, 65.79391, 66.24377, 66.32737, 65.94991,
    66.22871, 67.20421, 68.71222, 69.416, 70.12214, 70.8722, 71.48293,
    71.81638, 68.43542, 64.20288, 58.88104, 50.49883, 44.76797, 47.00963,
    44.16172, 42.3626,
  57.19136, 58.78287, 59.94012, 61.1394, 62.0788, 62.94897, 63.73335,
    64.42902, 65.05733, 65.61904, 66.13431, 66.58901, 67.01634, 67.28162,
    67.64862, 67.26617, 67.27358, 69.28852, 70.14197, 71.14231, 72.08765,
    72.85947, 73.3965, 73.73315, 73.61858, 66.45866, 48.74542, 44.69691,
    43.45109, 42.4829,
  57.43504, 58.88547, 60.03701, 61.16217, 62.09823, 62.97213, 63.71859,
    64.49635, 65.28973, 65.98164, 66.5257, 66.98185, 67.45441, 67.89473,
    68.30341, 68.54583, 68.83004, 68.35715, 69.22195, 70.84222, 71.98202,
    73.23518, 73.95423, 74.34882, 74.22578, 73.45561, 72.17574, 51.89093,
    43.58381, 42.37788,
  57.5667, 59.00539, 60.1864, 61.2238, 62.16336, 63.01897, 63.77556,
    64.44705, 65.22856, 65.90409, 66.58347, 67.49278, 68.1811, 68.54571,
    68.92947, 69.22828, 69.35648, 69.57031, 70.20111, 70.94323, 71.81709,
    72.48125, 64.04877, 67.9592, 68.34431, 73.85705, 73.68783, 72.95656,
    56.07211, 44.49989,
  57.89266, 59.20524, 60.44727, 61.43418, 62.2594, 63.15924, 64.00565,
    64.60256, 64.98976, 65.53805, 66.42785, 67.74153, 68.99626, 69.4966,
    69.82296, 70.16969, 70.22193, 70.24422, 70.68979, 71.31439, 71.53752,
    63.11929, 60.03945, 60.37749, 61.88797, 65.37718, 73.36662, 74.29774,
    74.19709, 54.54548,
  58.57531, 59.54602, 60.82867, 61.85499, 62.56999, 63.42478, 64.36011,
    65.12769, 65.51581, 65.82214, 66.42677, 67.5694, 69.08201, 69.70876,
    70.38546, 70.83599, 70.80435, 70.8834, 70.95036, 71.3247, 71.27921,
    60.19917, 64.15222, 63.24679, 62.66442, 62.44147, 64.37888, 73.47746,
    73.54919, 47.61771,
  60.82162, 60.69981, 61.67408, 62.37487, 63.08369, 63.8444, 64.69276,
    65.34654, 65.87537, 66.29984, 66.82442, 66.8815, 64.71111, 66.03111,
    66.75404, 67.61665, 69.55098, 69.25623, 67.57589, 67.25386, 64.89008,
    61.88572, 63.13682, 65.27874, 66.1354, 66.59661, 68.20434, 71.86763,
    64.67972, 41.37111,
  65.43172, 63.90834, 63.69763, 63.70138, 63.98537, 64.70593, 65.30292,
    64.37758, 64.06715, 64.58925, 65.06409, 64.38999, 64.6142, 65.19991,
    65.77971, 66.23515, 67.19904, 67.59642, 66.73698, 65.58414, 64.29527,
    63.35512, 63.05638, 64.26679, 66.42484, 71.63651, 73.68052, 70.03735,
    54.48609, 41.68461,
  71.37319, 70.12804, 68.03575, 66.65798, 66.01305, 65.85067, 64.71651,
    64.8811, 65.08147, 65.20453, 65.41763, 65.76562, 65.76314, 66.51056,
    67.10896, 65.62007, 66.32049, 68.24788, 69.56851, 68.90262, 67.8681,
    66.78526, 65.94528, 64.43681, 64.65063, 72.15794, 73.54716, 66.40529,
    41.60787, 42.10405,
  74.42345, 76.08768, 74.64059, 72.4071, 70.20381, 68.17756, 65.91481,
    65.99118, 66.02316, 66.26031, 66.07841, 66.20184, 66.47134, 65.60257,
    64.03027, 63.38287, 62.94884, 63.63034, 65.18637, 66.25355, 67.92723,
    68.23054, 68.31409, 67.897, 68.52077, 69.7748, 66.39113, 48.16521,
    41.77625, 41.61447,
  71.89853, 74.94946, 78.4595, 78.43956, 76.44393, 72.18857, 69.2998,
    67.84578, 67.1227, 67.67991, 67.0711, 66.41112, 66.48226, 66.76098,
    63.81535, 63.77657, 61.74752, 59.88099, 59.32006, 60.26296, 62.81129,
    63.62856, 64.67942, 71.47057, 73.03619, 72.61919, 52.20041, 42.87479,
    42.88554, 41.75462,
  67.37659, 67.49395, 73.61975, 78.0419, 80.05556, 76.71751, 71.99891,
    68.81842, 68.30156, 68.10367, 67.85619, 67.44466, 67.82908, 67.90753,
    67.68327, 67.3027, 68.2176, 65.10686, 61.41791, 59.01642, 60.46621,
    60.45186, 58.31445, 62.98344, 70.91687, 66.74754, 42.08776, 47.5617,
    43.61114, 42.39885,
  61.52374, 63.08232, 65.00574, 68.83544, 73.09928, 75.29381, 70.65454,
    67.42939, 70.37405, 69.4792, 69.51847, 69.1529, 69.4536, 69.62411,
    69.22424, 68.00243, 68.74197, 69.72677, 70.38264, 64.54491, 63.61198,
    63.03926, 58.71324, 51.98782, 49.64882, 51.19445, 42.46814, 43.9758,
    44.13094, 43.04866,
  61.54984, 62.3951, 62.41895, 59.85958, 59.73426, 64.24432, 66.85441,
    68.84067, 67.97295, 69.26004, 70.14898, 70.52306, 70.62637, 70.69415,
    70.17113, 69.186, 68.74558, 69.59046, 70.6428, 70.61633, 65.55364,
    61.43578, 52.22851, 46.89717, 42.69932, 42.3468, 42.42887, 41.69602,
    41.93272, 42.26522,
  61.59336, 59.03342, 63.07432, 63.67611, 64.49068, 64.93584, 65.78899,
    66.43694, 67.32394, 67.96706, 68.75983, 69.42103, 70.3297, 70.91056,
    70.70251, 70.5938, 69.80599, 69.22955, 65.5833, 61.96561, 53.60958,
    52.59071, 48.37562, 44.12713, 44.51305, 43.36158, 42.6717, 42.12754,
    41.73543, 41.69787,
  57.30674, 59.55312, 60.63129, 61.98455, 62.51134, 64.08234, 65.62138,
    66.10416, 66.55656, 67.15936, 68.04234, 69.03352, 70.14579, 71.30557,
    71.46176, 71.24905, 71.21687, 68.39464, 60.28446, 56.22333, 52.47236,
    50.07311, 46.67667, 44.42802, 43.80968, 43.19022, 42.52251, 42.09367,
    41.82431, 41.73971,
  61.53503, 60.76874, 61.76694, 62.65236, 62.90197, 62.84813, 63.40028,
    64.99519, 66.36166, 66.43117, 67.03191, 68.54183, 70.08546, 71.00593,
    71.5931, 72.30592, 72.85867, 72.9903, 67.72456, 61.16534, 53.94542,
    51.20427, 47.98092, 45.20926, 44.25926, 43.55778, 42.55824, 41.86354,
    41.61354, 41.64426,
  71.1787, 66.931, 64.04503, 63.90531, 65.05465, 65.0518, 65.34983, 65.51533,
    66.22161, 65.82088, 66.716, 68.06076, 69.25407, 69.8232, 70.39112,
    71.47374, 72.94682, 74.37029, 74.76719, 69.74658, 59.77152, 52.96036,
    49.13279, 46.76683, 44.70316, 43.84816, 42.97316, 41.74391, 41.56544,
    41.5427,
  80.80717, 76.07957, 69.46436, 63.86686, 66.63568, 66.60596, 66.86995,
    66.80286, 66.53704, 67.05283, 67.79362, 67.41797, 65.30679, 63.62354,
    62.08202, 62.80367, 66.544, 71.09409, 72.88763, 72.30107, 66.9184,
    57.88902, 51.05651, 48.94547, 46.11316, 44.62739, 43.5833, 42.05199,
    41.53796, 41.60875,
  79.85306, 76.41203, 70.08876, 65.70134, 68.11388, 68.59238, 69.19112,
    69.29582, 69.39301, 69.8018, 70.02223, 69.94688, 70.76602, 68.07655,
    64.89968, 62.95034, 62.54494, 63.5597, 63.98937, 63.72758, 62.79207,
    59.63628, 54.12427, 50.64339, 47.81808, 45.64495, 43.84739, 42.42498,
    41.50718, 41.65031,
  80.42207, 76.89757, 71.28495, 67.01505, 69.50893, 70.11008, 71.26965,
    72.14657, 73.11856, 72.95188, 71.73822, 70.32111, 71.15186, 71.10805,
    69.09954, 68.21651, 67.38051, 66.3987, 64.61466, 61.46181, 59.13583,
    58.15023, 56.07136, 52.18023, 49.61235, 46.4534, 44.46038, 42.46085,
    41.5542, 41.60968,
  80.53474, 77.52758, 71.34881, 67.90035, 70.88133, 71.644, 73.19218,
    74.12668, 75.82713, 77.17681, 76.15277, 75.30692, 74.66355, 73.70274,
    72.46837, 71.29496, 70.2877, 68.83556, 66.93109, 63.22628, 59.58863,
    56.53178, 56.2134, 52.83424, 51.05183, 47.85685, 45.231, 43.3283, 41.891,
    41.58789,
  80.97196, 78.31245, 71.84189, 67.99944, 71.2162, 73.07123, 74.98047,
    75.92569, 77.53107, 79.07579, 80.34181, 81.17291, 81.63961, 81.39615,
    79.58108, 77.77464, 76.20648, 73.65672, 70.96113, 67.4319, 63.17579,
    59.09703, 56.57799, 53.26987, 52.01779, 49.55431, 46.37646, 44.36399,
    42.89755, 41.9696,
  81.43464, 78.22448, 72.06768, 68.46115, 70.21725, 71.36671, 73.79119,
    76.20334, 78.35342, 79.97504, 81.1873, 83.37589, 85.64234, 86.75859,
    85.86674, 84.75509, 82.40644, 79.37067, 76.24039, 72.83047, 69.34549,
    64.55969, 59.41628, 55.68787, 53.74036, 51.81201, 49.01045, 45.68894,
    44.0198, 42.87168,
  81.73175, 77.65912, 69.53526, 64.51597, 65.38419, 65.74854, 68.31231,
    71.70751, 76.00449, 76.67126, 76.97543, 79.45824, 83.05681, 84.71049,
    82.88916, 81.80582, 79.90762, 77.60121, 75.25381, 72.97931, 69.9646,
    65.99281, 60.68637, 56.64399, 54.69228, 52.47568, 50.50726, 46.72083,
    44.23257, 43.30114,
  82.04507, 74.807, 67.75529, 62.07197, 61.78297, 60.97763, 62.80921,
    66.11614, 68.71899, 68.90475, 70.87283, 74.20395, 77.52954, 77.86771,
    76.3384, 75.16567, 74.21798, 71.96416, 70.17319, 68.90742, 66.74996,
    64.26031, 60.21748, 56.74804, 55.46386, 53.30815, 51.55815, 48.22175,
    44.21177, 42.87218,
  75.71516, 71.04069, 63.51791, 58.97147, 59.11833, 57.01695, 57.38731,
    58.62796, 59.45454, 59.51006, 61.6252, 64.89349, 68.52168, 69.45742,
    67.85109, 67.23745, 65.9267, 64.7833, 63.95803, 63.43363, 62.08635,
    60.42645, 57.54251, 55.15241, 54.54399, 53.38837, 52.46019, 50.36396,
    46.00774, 42.74232,
  64.36176, 62.69037, 58.0149, 55.57467, 56.66197, 55.80622, 53.89284,
    53.1339, 52.62584, 52.30951, 52.95275, 54.78172, 57.2448, 58.53704,
    58.04044, 57.46028, 56.43414, 55.4668, 55.73844, 56.5435, 56.11952,
    54.87306, 52.50049, 50.93373, 51.23877, 50.79068, 49.69323, 48.90689,
    47.47617, 43.70496,
  47.97906, 49.20826, 50.32523, 51.02106, 52.03776, 53.25647, 51.52185,
    48.42033, 47.42646, 47.83694, 47.51975, 47.27011, 47.14971, 47.61214,
    47.29527, 47.1107, 46.58231, 46.11761, 45.63396, 45.81094, 46.29981,
    47.44219, 47.95538, 47.46789, 47.70459, 47.69312, 46.97175, 45.06816,
    44.03468, 43.23487,
  44.65822, 45.36457, 45.94006, 45.66249, 46.31582, 47.69379, 48.11906,
    46.15154, 44.66988, 44.98771, 45.20568, 45.4476, 45.25974, 44.89572,
    44.52416, 44.23336, 43.55712, 42.72466, 42.58743, 42.55811, 42.40594,
    43.06377, 44.07186, 44.76011, 44.68679, 44.80246, 44.61723, 43.50667,
    42.44718, 41.80997,
  60.81105, 61.48001, 61.70709, 62.0791, 62.09572, 61.91135, 61.25101,
    60.12283, 58.81181, 57.66246, 56.72791, 55.96503, 55.18209, 55.34117,
    56.20119, 57.37299, 58.62656, 59.64368, 59.52978, 58.15707, 55.48675,
    51.84248, 48.70555, 46.35494, 43.43135, 39.09444, 36.20355, 37.88225,
    35.41198, 33.88988,
  63.08293, 63.64746, 63.45939, 63.75494, 63.96572, 64.2594, 64.41656,
    64.07639, 63.21037, 61.97977, 60.38256, 58.7311, 57.25744, 55.73362,
    54.70155, 54.88994, 56.20625, 58.85134, 61.93016, 64.49296, 66.14006,
    66.61884, 65.19398, 63.12344, 59.52267, 48.08649, 37.38216, 35.72523,
    34.94019, 34.08903,
  63.84554, 64.77986, 64.73688, 64.49571, 64.01003, 63.87152, 64.06654,
    64.54808, 64.96774, 64.90047, 64.03509, 62.72022, 61.00081, 59.31351,
    57.57017, 55.1383, 53.55283, 53.68556, 55.69151, 59.53239, 65.53233,
    71.1999, 72.60548, 70.53786, 66.31345, 60.74923, 54.71114, 39.37729,
    34.57791, 34.06932,
  64.72667, 65.68102, 66.43602, 66.93939, 66.81549, 66.41808, 65.66079,
    64.93372, 65.10422, 65.94711, 66.79668, 67.67117, 66.65845, 64.51305,
    63.22531, 61.67773, 58.97234, 55.91919, 54.69911, 56.24065, 60.79192,
    59.93574, 52.17388, 55.64872, 55.96713, 63.83117, 66.7832, 58.76453,
    43.64042, 35.47661,
  66.52776, 66.21303, 66.64462, 67.37669, 68.24124, 69.54039, 70.00187,
    67.83098, 66.12527, 65.29037, 66.77393, 71.72949, 75.00008, 72.93257,
    71.20441, 69.23492, 67.16936, 65.73748, 63.52905, 59.4917, 54.91459,
    49.28189, 45.93854, 47.7057, 49.72002, 52.74359, 60.59577, 73.53465,
    69.01015, 44.52623,
  68.41724, 68.78304, 68.44426, 68.05971, 68.3852, 70.96938, 71.95103,
    72.52512, 72.69547, 72.79897, 71.15433, 74.3125, 75.50356, 75.62989,
    75.92522, 73.19913, 67.99432, 70.12393, 72.34991, 66.03761, 57.57685,
    46.29055, 49.76633, 48.79074, 48.45545, 47.99138, 48.34051, 56.26642,
    60.22574, 39.25856,
  69.14629, 69.11067, 69.55035, 69.82278, 70.27147, 71.11397, 72.10336,
    72.77777, 73.24362, 73.54309, 73.84603, 68.81678, 56.31807, 56.3051,
    54.84534, 53.83107, 55.49024, 54.66177, 51.98735, 51.68205, 49.42646,
    47.85219, 49.72219, 51.85501, 52.31803, 51.69197, 52.03532, 54.94816,
    50.2074, 33.10684,
  71.43266, 70.37292, 70.31183, 70.40794, 70.75564, 71.57851, 72.0893,
    62.68388, 55.86422, 57.22707, 56.34526, 55.32193, 55.23943, 55.48936,
    55.71196, 55.38116, 54.59299, 53.3176, 51.52622, 49.80311, 48.3234,
    47.90812, 48.71907, 50.84949, 53.27011, 57.19537, 59.33455, 55.01968,
    45.36222, 33.3431,
  76.04851, 74.14411, 72.69954, 72.00867, 71.97298, 72.00811, 68.14602,
    63.84595, 60.74096, 57.56513, 55.9098, 54.64717, 53.95125, 54.91197,
    55.86312, 55.00059, 55.60255, 56.63907, 56.6892, 54.92899, 52.98219,
    51.61044, 50.56318, 49.17331, 50.48811, 57.93643, 64.09778, 53.93339,
    33.37505, 33.74446,
  81.22099, 80.32231, 78.10299, 76.0873, 74.82395, 73.40552, 71.57158,
    71.92597, 68.99549, 64.20507, 58.49273, 55.63303, 53.26956, 51.33343,
    50.02476, 50.33901, 51.07113, 52.23045, 53.70197, 54.70549, 55.80705,
    54.94704, 53.69668, 52.27752, 52.25796, 53.37585, 51.74184, 39.08471,
    33.37518, 33.34674,
  83.06567, 83.7336, 84.87716, 82.60917, 80.47371, 76.8137, 74.58932,
    73.28876, 72.84894, 73.68039, 66.57838, 58.1284, 54.50524, 50.74875,
    47.99158, 47.18963, 46.11664, 45.68251, 46.41408, 48.20371, 51.14912,
    51.86941, 52.06121, 57.51028, 65.44066, 61.64544, 42.28561, 33.85981,
    34.45773, 33.4259,
  80.66854, 80.74052, 85.14873, 87.32887, 86.57542, 82.43086, 77.95214,
    74.52017, 73.36737, 73.56029, 73.31131, 70.20134, 66.83534, 61.80942,
    55.59882, 51.1625, 50.48219, 47.97353, 45.80353, 45.06547, 47.32577,
    48.2136, 46.64328, 49.25229, 56.08363, 54.1615, 33.94434, 38.38849,
    35.00381, 33.96599,
  72.27824, 74.13045, 76.59178, 80.04423, 83.11184, 83.61415, 77.82722,
    73.26653, 75.812, 74.59499, 74.50401, 74.07588, 74.44122, 74.66264,
    72.00329, 55.0088, 57.46009, 57.65516, 54.5079, 48.81998, 48.73306,
    49.4675, 47.17092, 42.08955, 40.7855, 42.18062, 34.34664, 35.91165,
    35.68874, 34.56357,
  69.44855, 65.65855, 62.21022, 60.66497, 61.64768, 69.3924, 74.27298,
    75.52621, 70.8327, 74.10538, 75.19549, 74.9094, 74.83302, 74.99274,
    74.11005, 64.46581, 60.62991, 64.75607, 67.33316, 57.96437, 50.51329,
    46.39429, 39.47116, 36.28529, 33.89993, 34.00955, 34.08426, 33.49553,
    33.7792, 33.91865,
  67.56243, 63.01057, 64.28346, 62.82699, 62.14497, 61.89932, 63.07673,
    63.40977, 63.63564, 62.74342, 62.29898, 60.79554, 62.44307, 63.20432,
    64.70429, 70.44604, 62.61839, 56.43462, 53.01512, 48.40551, 40.4279,
    40.36654, 37.89132, 34.64394, 35.38647, 34.90296, 34.34663, 33.79744,
    33.4421, 33.38559,
  59.37522, 61.21423, 61.56643, 61.9069, 61.63744, 62.40348, 63.37095,
    64.0926, 63.33412, 62.03183, 61.68204, 61.52335, 62.014, 63.10351,
    59.84756, 57.81413, 57.9288, 51.59629, 46.12564, 43.30764, 40.39405,
    38.47223, 35.99946, 34.90058, 34.93696, 34.81673, 34.23865, 33.76187,
    33.5065, 33.44202,
  61.81033, 60.7384, 60.56953, 60.55666, 59.90712, 59.1162, 59.31642,
    60.64806, 61.29221, 60.55532, 60.21642, 62.85926, 66.26551, 66.73491,
    63.90114, 61.99446, 59.05238, 55.57401, 50.3885, 45.89104, 41.10928,
    39.49214, 36.95037, 35.43625, 35.38208, 35.02528, 34.14571, 33.53746,
    33.34239, 33.36616,
  69.88961, 66.0058, 62.67087, 61.71655, 61.24926, 60.26958, 59.86985,
    59.62875, 59.43753, 58.09459, 58.37689, 59.09547, 60.10682, 61.42297,
    61.33012, 62.98964, 63.79808, 62.39409, 58.98643, 53.38138, 45.49585,
    40.61455, 37.89784, 36.61444, 35.72968, 35.24229, 34.41845, 33.45604,
    33.32414, 33.31957,
  85.29389, 77.44703, 67.3513, 61.76098, 62.79877, 61.79364, 61.34597,
    60.67628, 59.24158, 58.50852, 58.02343, 56.19427, 52.8235, 51.11988,
    50.07567, 51.42268, 55.51768, 59.94946, 60.72571, 58.81436, 52.59061,
    44.78617, 39.76927, 38.52523, 37.00383, 35.99227, 34.98046, 33.67931,
    33.27951, 33.3331,
  83.30833, 77.38049, 68.37991, 63.37309, 64.2354, 63.54068, 63.19963,
    62.41432, 61.77055, 61.46789, 60.6734, 59.04097, 57.69718, 53.48542,
    49.728, 47.55978, 47.59094, 49.49272, 50.84834, 50.86793, 49.84074,
    46.65588, 42.24575, 40.03131, 38.21843, 36.65216, 35.22504, 33.94629,
    33.26953, 33.37048,
  81.93745, 77.22166, 68.38408, 64.23609, 65.27954, 64.87466, 64.91592,
    64.73104, 64.47405, 63.59828, 61.68596, 59.67238, 59.04578, 57.49562,
    54.63333, 52.64861, 51.08822, 49.86946, 48.39256, 46.29346, 45.21067,
    45.35728, 44.05268, 41.3194, 39.59101, 37.23607, 35.68873, 33.98995,
    33.30695, 33.37125,
  79.29462, 75.90506, 67.24641, 63.69077, 65.49936, 65.35449, 65.93892,
    66.39301, 67.0451, 66.90261, 64.92595, 63.25628, 61.65579, 59.77199,
    58.06097, 56.43062, 54.49913, 52.81076, 50.66623, 46.84329, 43.64857,
    42.64893, 44.53014, 41.81384, 41.0394, 38.5941, 36.41716, 34.65231,
    33.50393, 33.3288,
  75.69704, 73.24992, 65.08836, 61.71091, 64.17587, 65.18027, 66.0784,
    66.67778, 68.24986, 69.22799, 68.91823, 68.74684, 68.34085, 66.95512,
    64.82047, 62.89674, 61.01, 58.48433, 55.53617, 51.84305, 47.30435,
    44.47469, 44.4317, 42.19763, 42.14748, 40.24915, 37.61794, 35.68452,
    34.32273, 33.57349,
  72.12471, 69.24024, 62.64874, 60.12709, 61.7162, 62.33891, 63.96779,
    66.11794, 69.26346, 70.92576, 71.02663, 73.49869, 74.84624, 75.38065,
    73.25022, 71.47617, 68.69099, 65.71847, 62.035, 57.90398, 54.40012,
    50.75969, 46.47583, 44.30166, 43.62523, 42.31722, 39.76556, 36.8319,
    35.36204, 34.2908,
  69.8253, 65.21791, 58.78849, 55.42583, 56.34405, 56.82671, 59.35302,
    62.94432, 67.26094, 67.91031, 67.91596, 69.95328, 72.77332, 73.37447,
    71.75901, 70.68372, 68.72129, 65.99889, 63.40437, 60.41663, 56.56299,
    52.53059, 48.11636, 45.53309, 44.45974, 42.59934, 40.82449, 37.5931,
    35.41573, 34.58066,
  69.22438, 63.71735, 57.48314, 53.32128, 53.21286, 52.84108, 55.10402,
    58.8891, 61.75425, 62.08339, 63.75217, 66.29158, 69.05779, 69.11273,
    67.2104, 66.12785, 64.83112, 62.20474, 60.75483, 58.95499, 56.07697,
    52.93161, 49.21132, 46.75895, 45.92799, 43.46842, 41.55487, 38.46261,
    35.14301, 34.17799,
  65.48717, 60.81799, 54.70826, 50.66368, 50.72253, 49.42007, 50.25209,
    51.87764, 53.29946, 53.77277, 56.03255, 58.76321, 61.55748, 62.33627,
    60.39098, 59.60848, 58.26509, 56.96216, 55.67016, 55.569, 53.00291,
    50.91557, 48.30572, 46.5601, 45.9212, 44.33409, 42.93191, 40.62088,
    36.61155, 34.17282,
  56.32261, 54.27291, 49.67431, 47.18137, 47.82301, 47.62674, 46.79539,
    46.23986, 45.59803, 45.63825, 46.32507, 47.99232, 50.19475, 51.17063,
    50.85673, 50.22603, 49.53222, 48.37257, 48.95508, 49.39791, 48.45961,
    46.47866, 44.18491, 43.01226, 43.06035, 42.01897, 40.73139, 39.88277,
    38.31124, 34.96486,
  40.68272, 41.44444, 42.15465, 42.49164, 43.30755, 44.70605, 43.3417,
    40.371, 39.48841, 39.65377, 39.38542, 39.05128, 39.05083, 39.57756,
    39.35473, 39.36454, 39.01088, 38.59789, 37.98677, 38.19951, 38.6842,
    39.4674, 39.68537, 39.32931, 39.41924, 39.00967, 38.00847, 36.49054,
    35.6191, 34.75733,
  36.87737, 37.32011, 37.77193, 37.65869, 38.06649, 39.40715, 39.76044,
    37.5926, 36.43163, 36.7193, 36.94674, 37.23792, 36.93301, 36.58596,
    36.31836, 36.02529, 35.37285, 34.621, 34.47412, 34.46725, 34.3721,
    35.04738, 35.93472, 36.50143, 36.5477, 36.52969, 36.061, 34.97501,
    34.14098, 33.52433,
  49.95163, 49.76555, 49.3109, 48.73795, 47.97124, 47.16333, 46.39208,
    45.74042, 45.33132, 45.32843, 45.95731, 46.71184, 46.96366, 47.82017,
    48.46999, 48.54268, 48.13182, 47.32579, 45.73092, 43.68908, 41.22324,
    38.45515, 36.95572, 36.7057, 35.76355, 32.54873, 30.33326, 31.88206,
    28.27987, 26.8506,
  53.26037, 53.25456, 52.74205, 52.50912, 51.87652, 51.19089, 50.48459,
    49.57204, 48.56837, 47.58021, 46.99739, 47.18804, 47.79185, 48.16148,
    48.89587, 50.35071, 51.91983, 53.81143, 55.22261, 56.05053, 55.88747,
    54.62906, 52.49825, 52.02987, 52.10723, 42.15616, 28.82492, 30.22978,
    28.12767, 27.06895,
  54.35879, 54.55609, 54.15421, 53.85922, 53.48479, 53.32558, 53.33504,
    53.35556, 53.02938, 52.28131, 51.07402, 49.73652, 48.556, 47.72313,
    47.06812, 46.31042, 47.10411, 49.51608, 52.7877, 56.93287, 63.01768,
    68.57046, 68.18404, 64.5066, 60.03329, 51.77132, 41.62108, 31.37109,
    27.52276, 27.10806,
  55.69807, 56.55415, 56.67693, 56.69271, 56.30449, 55.99924, 55.69091,
    55.60904, 55.97123, 56.41354, 56.94148, 57.41322, 56.13275, 53.88505,
    52.59908, 50.83351, 48.46465, 47.5498, 49.78344, 53.50311, 58.55751,
    58.31026, 54.07813, 57.66767, 55.01655, 54.20054, 54.3323, 45.16648,
    33.09591, 27.77614,
  55.46298, 56.81166, 57.82401, 58.61701, 58.59068, 58.69903, 58.6785,
    57.11207, 56.18259, 56.18046, 58.17056, 63.76714, 67.49472, 65.86733,
    65.39584, 64.57575, 60.85396, 56.14927, 55.00069, 56.67861, 52.86875,
    42.52329, 42.95832, 47.02122, 51.20553, 54.33029, 58.71598, 65.82681,
    57.3343, 35.42329,
  54.61057, 55.93079, 57.48281, 59.13255, 59.74673, 62.00828, 66.61688,
    67.43516, 64.98401, 62.21411, 62.21113, 67.90894, 75.31764, 73.29961,
    74.43616, 75.69557, 72.73804, 67.64751, 62.14103, 57.83464, 49.70152,
    39.66747, 43.16161, 44.22459, 46.90998, 50.47738, 56.22145, 66.67161,
    59.63358, 30.12747,
  55.95513, 55.90508, 56.79829, 58.00302, 59.26257, 63.06631, 70.8097,
    76.48804, 77.17729, 73.04683, 68.5929, 59.38511, 47.81488, 48.04059,
    47.68465, 47.9618, 49.14768, 47.43893, 46.22328, 46.73699, 44.62592,
    42.86251, 44.13398, 45.91331, 46.75592, 47.63989, 52.22607, 57.08493,
    45.11172, 26.11065,
  61.94807, 59.84006, 59.51254, 59.42212, 60.1961, 64.95005, 66.89764,
    53.82481, 48.96875, 51.05071, 50.31642, 49.09137, 48.59837, 48.39408,
    48.06794, 47.73769, 47.27002, 46.05739, 44.31697, 43.66581, 43.89526,
    44.66068, 46.16933, 47.83587, 48.74992, 51.80556, 57.26499, 54.31986,
    37.40211, 26.34432,
  74.90125, 70.44473, 66.86767, 65.42577, 66.00085, 63.54438, 49.73538,
    47.72005, 48.00352, 47.69383, 48.192, 48.59111, 49.20319, 51.34171,
    52.68498, 51.26783, 51.58399, 52.03965, 51.33925, 48.90697, 46.83293,
    47.05228, 48.27233, 48.71257, 50.40232, 56.02223, 57.24866, 46.12937,
    26.59889, 26.82232,
  80.46468, 80.06738, 78.91502, 77.62991, 77.0661, 68.08478, 50.93441,
    52.95132, 49.58411, 47.28666, 45.58393, 46.10081, 45.76197, 45.07119,
    44.873, 46.97548, 48.86155, 50.15448, 51.06865, 51.79284, 52.31023,
    50.06122, 48.28053, 47.2365, 52.57788, 59.08222, 50.39016, 32.35536,
    26.39776, 26.21137,
  84.66625, 84.31385, 85.28344, 82.73544, 81.4508, 76.46256, 65.20895,
    62.37876, 59.02375, 55.2243, 47.15743, 41.98042, 41.34574, 39.91684,
    38.98888, 39.20878, 39.64151, 40.37751, 42.08334, 45.09194, 49.5185,
    49.9769, 48.31796, 51.67014, 56.10852, 51.28136, 35.02014, 26.69098,
    27.43725, 26.29073,
  87.87164, 87.35512, 90.00803, 90.61884, 87.74525, 83.43546, 79.4368,
    70.51544, 65.23278, 60.71011, 55.81501, 52.25806, 49.55285, 47.79007,
    45.43803, 41.74555, 41.35913, 39.87998, 38.91778, 39.61256, 43.36139,
    45.37337, 45.16643, 51.8354, 56.71048, 45.48677, 27.09844, 31.15382,
    28.0222, 26.86544,
  79.44205, 81.65994, 84.11671, 86.42556, 87.75001, 86.28169, 79.1562,
    73.28133, 76.31937, 70.36366, 64.61661, 61.73854, 60.78585, 61.90807,
    60.26684, 46.57388, 48.96341, 48.55799, 46.10854, 42.35327, 43.10646,
    43.75357, 40.84448, 36.63281, 36.41403, 34.92125, 27.77935, 29.34445,
    28.89748, 27.52992,
  59.36878, 56.67598, 55.13041, 54.3136, 55.72956, 61.25848, 68.81447,
    71.54642, 58.88183, 61.78247, 65.93314, 62.49934, 59.84071, 61.14919,
    60.09032, 55.46196, 54.2349, 57.9427, 61.08391, 52.7839, 46.31601,
    42.42567, 35.65156, 29.81943, 26.95687, 27.39653, 27.0342, 26.64886,
    26.98954, 26.94205,
  59.16158, 55.37618, 55.67475, 53.93358, 52.69732, 51.88315, 52.78173,
    52.95255, 50.91092, 50.21311, 49.7638, 48.92632, 51.32489, 51.4406,
    54.25248, 61.57814, 53.61289, 50.03535, 48.33291, 44.92903, 37.1986,
    34.64095, 30.0846, 28.04673, 28.54684, 27.92296, 27.34586, 26.8286,
    26.46837, 26.35558,
  50.61405, 53.07259, 54.06239, 54.68362, 55.06691, 56.35234, 57.49731,
    57.14822, 54.53596, 51.53976, 50.4529, 48.99519, 48.76029, 50.22218,
    47.76167, 46.6783, 47.51715, 42.33735, 38.27919, 35.38774, 32.12615,
    31.19128, 28.98259, 27.96796, 28.00333, 27.84344, 27.208, 26.85379,
    26.58179, 26.42156,
  49.21074, 48.18581, 48.31223, 48.86118, 49.38536, 50.07963, 51.59601,
    53.85554, 54.88838, 53.96792, 52.5433, 54.63522, 57.54387, 56.38419,
    51.8917, 49.75094, 47.03898, 44.53487, 41.2207, 37.58702, 32.78654,
    31.79745, 29.61188, 28.26357, 27.98674, 27.75558, 27.05681, 26.46324,
    26.34674, 26.30667,
  55.37844, 51.86563, 48.83851, 47.8937, 47.67577, 47.54417, 48.08796,
    49.37492, 50.55307, 50.72969, 52.79052, 54.78697, 55.6847, 56.40212,
    55.07654, 55.14551, 54.7262, 53.01273, 49.64376, 43.8497, 36.10722,
    32.6142, 30.42284, 29.341, 28.32403, 27.73998, 27.16459, 26.36934,
    26.25494, 26.23246,
  70.77393, 62.89122, 53.55347, 47.8679, 48.43822, 47.3189, 47.14737,
    46.97831, 46.32473, 46.49154, 47.2336, 46.5735, 44.47917, 44.67327,
    44.90255, 46.84577, 51.18552, 55.11042, 54.62555, 50.82257, 43.37619,
    36.16993, 32.03824, 30.87431, 29.39108, 28.44556, 27.6223, 26.57263,
    26.2315, 26.26416,
  71.34062, 64.77726, 56.20655, 50.59145, 50.97281, 49.98924, 49.45969,
    48.91803, 48.7076, 48.90068, 48.18037, 46.06845, 45.39714, 42.66379,
    40.5037, 39.70272, 40.95548, 43.7556, 45.02905, 44.33331, 42.23844,
    38.53233, 34.56185, 32.44122, 30.74718, 29.08481, 28.02495, 26.74303,
    26.21613, 26.27261,
  72.49151, 67.26952, 58.95329, 54.13097, 54.29472, 53.34652, 53.02886,
    52.53254, 52.04393, 51.26955, 48.99294, 46.95773, 47.18118, 45.85714,
    44.05385, 43.02217, 42.63657, 42.65074, 42.27034, 40.29311, 38.77706,
    38.15933, 36.39148, 34.08375, 32.06671, 29.78166, 28.18888, 26.79559,
    26.22799, 26.2598,
  72.45596, 69.00632, 61.02569, 57.39697, 58.30231, 57.43313, 57.37735,
    57.19859, 57.22671, 56.17043, 53.3553, 50.98729, 49.632, 47.87209,
    46.13221, 45.02844, 43.96082, 43.40788, 42.76806, 41.39305, 39.65063,
    37.69898, 36.48148, 35.41562, 33.78759, 31.00926, 28.80601, 27.33182,
    26.35365, 26.23884,
  70.62356, 68.2489, 60.94695, 57.83809, 59.83935, 60.32595, 60.48499,
    60.44975, 61.38444, 61.28706, 59.8868, 59.31778, 58.05698, 56.02108,
    53.39021, 51.24586, 48.96156, 46.50367, 44.47746, 42.36074, 40.42525,
    38.15387, 36.11879, 35.44423, 35.42385, 32.94904, 29.98825, 28.2785,
    27.14164, 26.39282,
  67.13259, 64.75594, 58.8855, 56.59, 57.69377, 57.84418, 58.97409, 60.81722,
    64.2459, 64.97128, 64.12568, 66.29221, 67.20117, 67.05761, 64.25288,
    61.64311, 58.20359, 54.32014, 50.443, 46.661, 43.67766, 40.98593,
    38.29848, 36.64568, 36.42471, 35.48649, 32.82418, 29.57073, 28.24869,
    27.06288,
  64.77299, 60.49578, 54.47263, 51.18151, 51.57766, 51.76742, 54.1754,
    58.24129, 63.03073, 62.76304, 61.7692, 63.81411, 65.88442, 65.83816,
    64.17294, 62.55347, 59.69743, 56.45087, 53.50584, 50.516, 46.38424,
    42.92731, 39.56137, 37.38324, 37.01139, 36.08076, 34.5974, 31.05996,
    28.64247, 27.56291,
  62.72053, 58.41183, 53.20081, 49.07102, 48.46692, 48.05895, 50.7949,
    55.2369, 58.41236, 57.90922, 59.18954, 61.2822, 63.28864, 62.68498,
    60.57006, 59.90585, 57.71999, 55.22887, 53.51154, 51.41137, 48.05547,
    44.80383, 41.54866, 39.49076, 38.81369, 37.33479, 35.76026, 32.17849,
    28.20552, 27.07425,
  59.29367, 55.15868, 50.06757, 46.51971, 46.33713, 45.02347, 46.38868,
    48.69052, 50.23448, 50.691, 52.4282, 55.04356, 57.38997, 57.43503,
    56.42519, 55.52226, 53.73353, 51.42556, 50.55807, 49.40716, 46.42591,
    44.43871, 42.23739, 40.51728, 40.09032, 39.18311, 38.32127, 35.3998,
    29.83463, 26.88525,
  52.55026, 49.9053, 46.15216, 43.76685, 44.34946, 43.89791, 43.15721,
    42.50473, 41.68456, 42.00257, 42.80107, 44.52754, 46.68747, 47.50162,
    47.27553, 47.00569, 45.76487, 44.53921, 44.64954, 44.58282, 42.81351,
    40.1009, 37.41177, 36.30045, 36.56761, 36.11264, 35.41337, 34.81103,
    32.57635, 28.12632,
  37.14623, 37.81565, 38.23145, 38.40808, 39.37299, 40.80145, 38.87083,
    35.51556, 34.54134, 34.97304, 34.85785, 34.69359, 34.7718, 35.00852,
    34.7898, 34.57608, 34.27036, 33.66002, 32.95172, 33.00256, 33.15255,
    33.40695, 33.03075, 32.27689, 32.45803, 32.34852, 31.58087, 29.97226,
    29.19567, 28.08179,
  31.78664, 32.42253, 32.66209, 32.1549, 32.50372, 34.25742, 34.90364,
    31.72127, 30.33959, 31.06425, 31.59221, 32.03507, 31.90606, 31.35583,
    30.77664, 30.35084, 29.18088, 28.17638, 28.00438, 27.93086, 27.8356,
    28.4297, 29.15909, 29.61448, 29.74265, 29.79848, 29.342, 28.15177,
    27.0956, 26.35501,
  41.0709, 40.70198, 40.56442, 40.59738, 40.59343, 40.89241, 41.39704,
    41.99414, 42.74264, 43.73611, 45.22152, 45.75439, 44.28613, 44.66003,
    45.07596, 44.9068, 45.16792, 45.99405, 46.72889, 47.37283, 46.95552,
    45.22814, 45.1007, 46.33414, 46.76379, 44.98433, 45.43275, 46.7686,
    38.31458, 35.5373,
  44.52048, 44.22018, 43.39281, 43.32419, 42.64465, 42.22436, 42.40002,
    42.8248, 43.57603, 44.73753, 46.43492, 48.72148, 50.67912, 50.92096,
    51.54832, 53.23882, 54.21434, 56.33661, 58.43306, 60.01078, 59.86456,
    58.6074, 57.51735, 58.80151, 60.0772, 51.96653, 42.22549, 44.61995,
    38.43477, 36.30056,
  46.52267, 46.90657, 47.00663, 46.94008, 46.74759, 46.46882, 45.96954,
    45.62069, 45.5014, 45.53749, 45.85554, 46.86898, 48.43126, 50.67667,
    52.77926, 53.2726, 55.44049, 58.875, 62.45352, 66.99094, 72.92011,
    74.39527, 74.42875, 74.44418, 70.01521, 61.47487, 52.49731, 44.4276,
    37.86341, 36.70858,
  49.03335, 49.61426, 50.42759, 51.22614, 52.0123, 52.86174, 52.91119,
    52.5828, 52.69449, 52.74918, 52.7552, 53.06177, 52.69348, 52.05466,
    54.07308, 55.57656, 54.47294, 54.14654, 58.57062, 64.42964, 71.39616,
    72.0529, 68.74593, 72.33113, 69.28313, 66.23376, 62.31182, 52.72575,
    41.64776, 36.38276,
  51.689, 51.90981, 52.83856, 53.33118, 53.66866, 54.10713, 54.71555,
    54.92451, 56.19132, 57.48702, 58.90456, 63.36036, 66.21749, 65.49455,
    66.06325, 66.6772, 63.78055, 59.23833, 59.90742, 64.81767, 64.06285,
    56.54979, 58.10656, 63.74734, 68.32693, 68.70875, 66.78141, 71.04931,
    64.10095, 43.46228,
  51.92118, 54.2637, 56.22755, 58.01376, 57.56094, 58.35981, 62.09696,
    62.80856, 61.86579, 61.43927, 63.88245, 70.12928, 71.17995, 71.42616,
    72.37431, 73.4012, 73.16143, 72.20278, 67.4846, 65.72792, 59.79349,
    52.35574, 56.92306, 60.19492, 64.2466, 65.58176, 66.65398, 73.78519,
    67.45148, 39.10558,
  49.71597, 52.89402, 55.97879, 58.9879, 60.35203, 63.5827, 70.58958, 71.28,
    70.77723, 70.27016, 67.38636, 60.06591, 50.99709, 53.27687, 55.76213,
    58.33406, 60.00471, 58.32607, 55.43526, 57.2681, 56.13543, 55.92011,
    58.87757, 62.60412, 63.14013, 60.85051, 63.91162, 67.6202, 55.81628,
    34.76509,
  49.57835, 51.40582, 54.93132, 58.44321, 61.11434, 67.53252, 71.02744,
    59.87332, 55.07638, 57.13472, 56.3176, 55.20993, 54.92492, 56.52559,
    57.54272, 58.54747, 60.26382, 59.87821, 57.33667, 57.22947, 58.04506,
    60.74501, 64.55499, 66.57884, 64.756, 65.74364, 70.71736, 66.46037,
    49.64321, 35.32675,
  63.65012, 60.84318, 59.88868, 60.53326, 61.17865, 61.61034, 53.66201,
    54.48262, 57.83565, 60.10639, 62.03503, 63.12587, 64.63702, 70.54762,
    73.84943, 67.95212, 68.53681, 70.94675, 70.59913, 66.10562, 63.06762,
    66.26547, 70.75852, 70.24332, 67.14542, 72.84898, 72.25103, 58.57199,
    36.87547, 35.75789,
  74.99737, 75.53878, 74.26521, 73.50508, 72.0062, 64.61495, 50.07636,
    54.70578, 54.30121, 56.21215, 58.63419, 62.37751, 62.13873, 60.87293,
    60.04749, 64.84971, 67.88863, 69.21241, 69.76562, 71.92432, 73.6961,
    69.44364, 65.04034, 60.09601, 65.1562, 72.21693, 62.2215, 43.82201,
    35.27571, 34.12883,
  75.44606, 75.88941, 78.01404, 75.13, 74.41441, 72.60906, 64.50189,
    64.74209, 65.19623, 64.64053, 55.60518, 46.05655, 44.6072, 45.23552,
    45.95645, 48.00124, 50.22396, 51.94642, 54.35608, 59.88279, 69.24406,
    67.51156, 59.34645, 59.64841, 64.01814, 59.79525, 44.10563, 35.85909,
    36.10231, 34.34452,
  79.86385, 77.9912, 80.20001, 81.40247, 79.00703, 76.20745, 73.3951,
    70.28583, 63.16079, 60.52779, 57.18129, 54.28209, 55.93378, 54.56132,
    48.80974, 48.83044, 48.34644, 48.44629, 48.92113, 52.18872, 59.72398,
    62.13668, 56.36819, 63.18434, 65.79482, 53.62094, 36.14709, 40.19313,
    37.21508, 35.36499,
  78.09135, 79.50847, 81.03492, 82.63487, 82.77872, 80.58684, 73.47889,
    69.7449, 71.77466, 70.29989, 70.53113, 70.21159, 71.30314, 71.94954,
    65.99145, 54.3954, 55.24902, 55.32305, 53.99853, 54.83013, 57.70335,
    56.95795, 52.29, 48.11083, 47.3339, 44.31703, 36.83023, 38.49717,
    38.35266, 36.3297,
  71.39421, 73.10712, 67.96981, 67.62688, 68.3788, 71.48201, 72.36886,
    72.67346, 70.9866, 72.04446, 72.8119, 72.18168, 73.25797, 73.4763,
    72.33137, 69.97717, 62.37225, 67.48561, 70.22437, 63.80914, 56.86314,
    52.55462, 46.01466, 40.37356, 37.44852, 37.07101, 35.92781, 35.41335,
    35.87518, 35.58027,
  59.10861, 57.28467, 59.21856, 59.35253, 60.93741, 66.23096, 72.85117,
    69.09874, 65.73772, 65.42233, 63.19411, 60.60003, 63.83717, 70.50945,
    71.69632, 68.25157, 64.05644, 62.29718, 63.50899, 59.32204, 47.39501,
    45.79897, 40.42935, 38.66259, 38.81018, 37.56055, 36.49083, 35.68365,
    35.03123, 34.67712,
  54.41165, 57.96643, 59.56352, 60.15263, 60.17997, 62.29035, 65.46375,
    64.58066, 59.73649, 56.66193, 56.53154, 54.5522, 53.681, 57.14425,
    55.40199, 55.17323, 57.13825, 53.51412, 52.13933, 48.50765, 41.6991,
    42.47352, 39.20271, 38.11004, 38.25262, 37.66937, 36.15022, 35.71506,
    35.24048, 34.76601,
  46.98098, 46.83472, 48.64312, 51.24928, 53.86547, 56.37258, 59.09414,
    62.71999, 64.2205, 62.63525, 59.28667, 63.25386, 69.33112, 65.91492,
    58.1972, 55.88013, 53.31438, 52.32042, 52.65342, 49.58516, 41.6809,
    42.9468, 40.21698, 38.5112, 37.83844, 37.53408, 35.88005, 34.70977,
    34.65069, 34.53902,
  46.55049, 45.19782, 43.67196, 44.9416, 46.68554, 48.99207, 51.73667,
    55.20176, 57.87569, 59.2317, 64.72781, 69.5183, 70.16285, 71.67419,
    68.01048, 65.23923, 62.79734, 62.13981, 61.24042, 54.72744, 43.78725,
    42.47046, 40.83185, 39.89289, 37.69281, 36.55339, 35.8978, 34.47023,
    34.41233, 34.31447,
  59.77509, 52.97569, 44.55647, 40.24794, 42.06574, 42.60262, 44.26804,
    46.16086, 47.38512, 50.04373, 53.86667, 53.89734, 50.92596, 54.33013,
    56.65652, 60.14145, 67.12523, 73.75174, 73.97292, 66.66968, 53.92508,
    46.37512, 42.38486, 40.79007, 38.42622, 36.81421, 35.91294, 34.75216,
    34.35253, 34.31028,
  59.22413, 53.19474, 45.78539, 40.48006, 41.46334, 41.71899, 42.67839,
    44.01783, 46.31466, 50.05751, 50.40122, 45.30107, 46.04281, 45.83323,
    45.65571, 46.28807, 50.06751, 56.11727, 60.5554, 61.42615, 57.62179,
    51.52942, 45.67869, 42.72353, 40.3564, 37.68147, 36.28058, 34.92657,
    34.3544, 34.33152,
  61.15903, 55.38147, 47.6408, 43.06343, 42.89337, 42.48197, 42.85592,
    43.75835, 45.66074, 47.37894, 44.71823, 41.44024, 44.37728, 44.38815,
    43.53086, 43.36605, 44.92289, 47.43808, 50.52499, 51.90753, 52.65117,
    53.30239, 50.50211, 46.0526, 42.27389, 38.61613, 36.45302, 35.09541,
    34.3558, 34.33347,
  65.28211, 60.73647, 53.29326, 49.93913, 50.04028, 48.48914, 48.2732,
    48.06247, 49.85641, 50.04718, 45.65086, 43.15282, 44.26383, 44.13044,
    43.51891, 43.68475, 43.89294, 44.95549, 46.86087, 48.39399, 49.83033,
    50.31524, 50.77462, 50.09996, 46.17124, 40.29876, 37.20055, 35.83702,
    34.54372, 34.28971,
  67.16878, 65.65404, 58.44949, 55.99321, 58.14861, 58.6675, 57.7319,
    55.62717, 56.24251, 55.08324, 51.33263, 52.19829, 52.51118, 52.14027,
    50.36048, 49.93909, 49.16993, 47.37524, 46.85669, 47.20023, 48.02732,
    48.20166, 47.68561, 48.3735, 49.09676, 44.25793, 39.13235, 37.49527,
    35.83999, 34.50772,
  67.03204, 64.99949, 60.68145, 59.24008, 59.87777, 59.56493, 60.83027,
    61.46786, 65.21009, 63.41169, 59.31343, 62.55365, 64.58508, 65.23721,
    63.04847, 61.24973, 59.36332, 56.58586, 53.07663, 51.30445, 50.76848,
    50.21234, 48.69682, 47.81687, 48.70808, 48.75418, 44.51906, 39.49314,
    37.77253, 35.58383,
  66.30157, 62.0524, 56.3001, 53.63621, 53.9875, 53.80454, 56.12629,
    60.93273, 66.90712, 63.71505, 59.39072, 62.80761, 65.23955, 65.82226,
    64.7327, 64.19572, 62.41767, 61.09284, 59.14765, 56.95301, 55.36814,
    53.61044, 50.77147, 48.58431, 48.71285, 49.31611, 48.35146, 42.88153,
    39.17503, 37.02882,
  66.66309, 63.76265, 58.72377, 53.86076, 51.84546, 51.23871, 55.34786,
    61.21564, 63.38269, 59.99362, 60.7639, 63.11721, 65.21345, 64.46812,
    62.23576, 62.06329, 62.07579, 61.98353, 62.02813, 61.33776, 60.53613,
    59.59608, 56.46728, 53.67382, 53.06488, 51.81674, 50.68057, 45.32223,
    37.75571, 35.96353,
  63.63333, 59.70186, 54.80236, 51.59694, 50.41882, 48.30479, 51.05843,
    53.70116, 53.9391, 53.60993, 56.67195, 59.40855, 61.09805, 60.88593,
    60.10001, 59.52385, 59.27419, 59.55482, 60.61075, 60.84231, 60.52498,
    61.75436, 61.52899, 59.63376, 59.25328, 58.35228, 58.27171, 53.47821,
    41.23442, 34.96592,
  56.77265, 55.27276, 53.34213, 52.91795, 53.93655, 52.27303, 51.09933,
    49.26467, 46.25348, 47.79507, 49.53366, 51.94913, 54.16576, 55.26546,
    55.71947, 55.48321, 54.13286, 54.4236, 56.54921, 58.01033, 56.0115,
    53.35126, 50.82565, 50.58939, 51.8153, 52.35512, 52.64288, 53.83924,
    49.38321, 38.21014,
  45.42715, 46.18675, 47.05994, 48.65059, 52.40113, 56.24994, 52.67149,
    45.48821, 43.61414, 45.19711, 45.22538, 45.73511, 46.55886, 47.46072,
    47.93455, 47.94643, 47.35315, 46.81612, 45.95404, 44.86103, 44.63564,
    44.58407, 43.09643, 42.18281, 43.2294, 44.05884, 43.62227, 41.7001,
    41.18621, 38.87498,
  41.68302, 42.2997, 42.68707, 42.36013, 44.46715, 49.50209, 51.35947,
    44.41739, 41.54109, 43.86012, 45.65528, 47.36722, 48.06783, 47.45197,
    46.20102, 45.01338, 41.70195, 38.68848, 38.55615, 38.16735, 37.28402,
    37.94423, 38.4709, 38.75706, 39.22205, 40.11906, 39.95484, 37.84874,
    35.76109, 34.34846,
  40.18649, 40.48781, 40.74615, 41.08526, 41.19059, 41.47139, 41.88833,
    42.39307, 42.92025, 43.80946, 45.7424, 45.67905, 42.2917, 42.57827,
    42.88939, 42.40937, 42.70087, 43.75299, 44.81457, 46.55736, 47.06219,
    45.38131, 46.07779, 48.65045, 50.57195, 50.21921, 54.99167, 56.9692,
    42.51632, 39.09628,
  42.93496, 43.60371, 43.16237, 44.13511, 43.88202, 43.77835, 44.39709,
    44.93245, 45.5782, 46.33793, 47.56509, 49.42292, 50.53206, 48.51603,
    47.2446, 48.11365, 47.3138, 48.53128, 50.38308, 51.685, 51.17831,
    50.28732, 50.46935, 53.89856, 57.15062, 53.07907, 50.49022, 54.82548,
    43.355, 40.29144,
  42.60379, 43.38723, 44.30963, 45.12542, 45.79379, 46.3412, 46.51107,
    46.89923, 47.35231, 47.95745, 48.63748, 49.90467, 51.41517, 53.47969,
    54.78685, 52.87199, 53.1886, 54.88746, 55.95197, 57.717, 60.89408,
    64.09148, 65.35661, 65.84671, 65.20429, 60.59856, 57.65643, 53.48627,
    43.07086, 41.39546,
  45.46835, 46.24192, 47.63899, 49.049, 50.74373, 52.50218, 52.62471,
    52.05023, 52.33825, 52.87205, 53.28811, 54.14401, 53.9441, 53.13735,
    56.471, 58.69583, 55.65657, 52.89746, 55.61003, 58.84655, 63.70295,
    64.74656, 63.69058, 68.50137, 68.84442, 66.9677, 61.56152, 52.81737,
    44.16642, 39.64215,
  47.98704, 47.83244, 49.70293, 51.14157, 52.55194, 53.19638, 53.20741,
    53.38531, 54.68252, 55.64918, 56.06194, 58.86186, 60.38108, 60.70966,
    61.83413, 63.27111, 61.04104, 55.63723, 56.31476, 60.82685, 60.38531,
    54.71687, 56.65988, 63.40927, 70.09345, 67.92764, 59.65313, 62.39139,
    59.79251, 44.81553,
  49.50779, 51.90623, 55.36622, 58.52894, 58.68139, 59.16002, 61.55196,
    62.04459, 61.35904, 62.00301, 64.37285, 69.72532, 75.2344, 73.29542,
    74.83, 77.77551, 77.70103, 71.0479, 61.77258, 62.48888, 58.04005,
    52.69329, 56.30472, 61.59932, 67.35926, 65.90386, 60.6372, 68.57724,
    64.67519, 43.29624,
  50.25443, 52.78637, 56.15762, 59.15482, 59.70557, 60.78596, 63.69291,
    66.08396, 65.69136, 64.71765, 64.06814, 60.68958, 56.28954, 58.94284,
    61.46267, 63.50697, 66.29507, 63.07121, 55.99383, 58.0766, 56.42956,
    56.03279, 59.41875, 65.60314, 66.50919, 59.8721, 60.09998, 63.86243,
    57.31219, 39.48132,
  50.81591, 53.13725, 56.77331, 59.92318, 60.27595, 64.32588, 67.68596,
    59.76229, 54.90767, 56.22153, 56.1986, 56.30251, 57.04904, 60.72014,
    63.76284, 66.13126, 69.24874, 68.39101, 62.68374, 61.42087, 60.78774,
    62.92822, 67.92811, 70.72303, 66.56559, 64.27529, 68.88274, 66.45387,
    54.61208, 40.0879,
  60.08979, 61.08802, 62.88537, 63.16914, 61.58746, 63.68853, 61.35508,
    62.00868, 65.96465, 68.78712, 70.32806, 71.89495, 75.4715, 82.37556,
    84.14858, 81.49577, 82.27402, 83.44904, 82.96042, 77.61071, 72.01012,
    77.0642, 82.07333, 80.88503, 71.53514, 76.9132, 75.61798, 63.65864,
    43.51115, 39.42085,
  78.97967, 80.73521, 80.4772, 80.93198, 79.07312, 76.1227, 63.33824,
    68.20181, 69.85194, 77.54649, 81.68353, 83.09363, 82.59476, 80.88708,
    74.09148, 80.70741, 81.91133, 82.27957, 82.29476, 83.39276, 84.17135,
    81.85502, 77.19621, 68.38316, 67.68436, 70.30101, 64.01891, 47.69297,
    39.20781, 36.86443,
  77.19295, 76.73196, 78.53589, 78.31448, 79.48312, 79, 73.33273, 75.88558,
    79.02646, 78.1898, 70.04823, 54.71823, 53.19867, 53.67969, 55.02024,
    57.09474, 60.55373, 63.29168, 67.38402, 71.75893, 77.8839, 74.72444,
    58.03397, 54.30634, 57.08432, 54.574, 45.09793, 39.42807, 38.81422,
    37.00167,
  82.73386, 80.48251, 83.90919, 84.41138, 82.25327, 80.19894, 73.87919,
    68.494, 61.79405, 56.46909, 53.68917, 51.92387, 54.35485, 56.14128,
    56.02771, 56.1044, 56.39422, 59.93592, 66.84452, 74.23416, 75.7059,
    68.11109, 54.90739, 61.00962, 62.05085, 50.75774, 39.69246, 41.71143,
    40.20705, 38.17159,
  86.42857, 88.46391, 90.46785, 90.52644, 89.51033, 85.94711, 77.87772,
    72.72367, 76.32785, 65.56985, 63.79964, 61.50194, 64.77151, 67.5927,
    65.01688, 57.92742, 59.92165, 62.13633, 68.58102, 79.47099, 75.50498,
    61.37811, 53.6352, 50.92104, 50.82079, 46.61842, 40.56466, 41.54433,
    41.68034, 39.26184,
  76.80555, 77.62281, 78.32401, 77.56332, 77.32806, 78.04962, 79.4532,
    79.73878, 76.94855, 77.02414, 77.65585, 76.07705, 77.38538, 78.1881,
    74.97504, 66.0384, 63.68483, 66.71248, 70.90422, 69.28294, 60.91251,
    54.67294, 50.63525, 45.09463, 42.46427, 41.63183, 39.54301, 38.87165,
    39.24909, 38.58396,
  64.62951, 64.34718, 67.86902, 71.14379, 73.21976, 75.10336, 79.53381,
    80.13012, 76.2589, 75.0513, 71.06403, 67.9022, 72.20859, 74.13731,
    72.14268, 72.7756, 69.68552, 70.06696, 74.70368, 71.37796, 50.9701,
    50.2248, 45.38928, 44.21599, 43.36284, 41.52322, 40.11353, 38.987,
    38.0896, 37.55373,
  64.88821, 67.36932, 69.63715, 69.08097, 67.95583, 72.69852, 78.581,
    76.47732, 69.72272, 66.81348, 67.94405, 63.93141, 61.94458, 67.52411,
    64.79467, 64.48283, 67.14339, 64.22003, 65.23803, 61.97453, 46.60239,
    47.85269, 44.50777, 44.28291, 44.11903, 41.56218, 39.61478, 38.9718,
    38.29358, 37.60176,
  57.76333, 56.19147, 58.26015, 60.16018, 61.51789, 63.86118, 67.79693,
    71.59305, 72.20412, 71.19055, 66.10123, 71.83424, 80.78844, 76.73508,
    65.48464, 63.97067, 61.536, 60.24462, 64.31268, 62.69196, 45.82421,
    48.22802, 45.45618, 44.29207, 43.12307, 41.20412, 39.19233, 37.71852,
    37.63183, 37.38667,
  53.60335, 54.90339, 55.23473, 58.16568, 61.07548, 64.2032, 65.5607,
    65.84108, 66.25123, 67.49848, 76.60731, 82.33573, 82.39737, 80.39282,
    78.13354, 71.85426, 63.90728, 62.26315, 67.71128, 62.35625, 46.90234,
    45.8847, 44.28127, 43.79269, 41.05857, 39.54411, 39.04258, 37.23398,
    37.23151, 37.07222,
  59.04679, 55.86102, 50.78004, 48.40009, 50.54607, 51.6894, 53.92182,
    56.32389, 57.0106, 61.08912, 68.42336, 68.7403, 61.08422, 63.62686,
    66.77401, 72.57965, 83.10152, 85.63683, 84.74483, 76.60106, 57.84986,
    48.90961, 44.96945, 43.56877, 40.76891, 39.07739, 38.52578, 37.525,
    37.18467, 37.04854,
  57.58954, 55.48539, 50.75446, 47.24871, 48.80872, 49.82249, 51.02136,
    52.69158, 56.24788, 63.72827, 66.17048, 57.79666, 57.34759, 56.95722,
    56.74003, 58.30253, 65.09877, 71.63783, 70.74014, 69.46758, 63.70766,
    54.92204, 47.66372, 45.20147, 42.9032, 39.79281, 38.57167, 37.64369,
    37.1718, 37.0588,
  54.7061, 53.07392, 48.56087, 46.15324, 46.67099, 47.35178, 48.38424,
    50.0513, 53.80865, 58.80151, 56.05991, 50.4374, 54.73549, 54.87063,
    53.6147, 52.09193, 53.08345, 54.43001, 55.63299, 56.08772, 56.89033,
    58.80946, 54.80533, 49.89125, 45.29015, 41.12476, 38.75307, 37.6876,
    37.19529, 37.09351,
  55.85629, 51.15801, 48.38898, 47.35653, 47.9133, 46.84957, 47.84614,
    48.88086, 53.61021, 56.02075, 49.26533, 45.17324, 48.09176, 49.29637,
    49.40972, 50.01448, 50.25117, 50.84037, 52.50843, 53.56158, 53.78134,
    54.54435, 56.71224, 56.27795, 50.31803, 42.7293, 39.1615, 38.35132,
    37.43033, 37.07991,
  59.2438, 57.66503, 51.72387, 51.65667, 54.73083, 56.32972, 55.9254,
    53.85233, 55.57528, 54.98923, 47.98412, 48.32604, 49.6226, 50.90789,
    50.59655, 51.90169, 52.39577, 50.24427, 49.47888, 49.3791, 49.03288,
    49.0652, 49.32734, 51.66383, 53.88758, 48.09347, 41.79217, 40.32242,
    38.9855, 37.29415,
  65.78283, 64.43739, 60.66309, 61.29814, 62.33784, 60.98297, 66.39139,
    67.35196, 65.8848, 62.81274, 54.76693, 57.13277, 58.47736, 58.62636,
    57.48779, 58.19843, 58.21616, 56.36901, 52.89579, 51.25109, 49.79183,
    48.85789, 48.34088, 48.14823, 50.73632, 54.01951, 49.59693, 42.53481,
    40.79141, 38.28455,
  64.77323, 62.25859, 56.03258, 53.88116, 55.83085, 56.44034, 57.28156,
    60.64562, 66.61515, 62.92009, 54.00472, 56.06601, 57.11615, 58.37505,
    59.11503, 61.04491, 61.46374, 61.53084, 58.79893, 54.68996, 52.98386,
    52.00207, 50.57072, 49.07688, 49.33397, 52.50475, 53.94817, 47.89067,
    43.96107, 40.67464,
  69.63799, 69.4631, 64.88113, 58.35333, 56.44276, 56.53519, 61.1483,
    66.26227, 65.05386, 59.98255, 58.29285, 58.62675, 59.95185, 59.51991,
    58.27324, 60.02347, 62.26063, 63.34303, 62.81022, 60.25355, 58.29794,
    57.29305, 54.32726, 51.29846, 51.46917, 52.42135, 54.49532, 50.25908,
    42.11915, 39.55329,
  70.45502, 67.88185, 62.17431, 57.87844, 57.19882, 55.20668, 59.94849,
    62.3339, 58.58847, 56.63464, 58.79574, 59.11042, 59.02508, 59.13016,
    59.78276, 61.06395, 63.12492, 65.54013, 66.60234, 65.58891, 65.24881,
    67.45475, 67.50823, 63.37506, 61.76251, 62.51315, 64.25197, 60.48528,
    45.57557, 37.67134,
  67.45963, 63.46689, 63.32705, 63.32774, 65.61718, 63.82706, 62.9211,
    59.41564, 53.16123, 55.02897, 56.2211, 56.91326, 57.2311, 58.08922,
    60.05193, 60.65286, 60.38612, 61.29101, 63.26704, 66.23734, 65.62228,
    62.43447, 60.52545, 60.44792, 60.99408, 60.66869, 60.08101, 63.60462,
    58.53045, 42.3639,
  56.69877, 57.3046, 59.3335, 60.89741, 66.08687, 71.23193, 67.93445,
    56.88038, 52.77383, 54.24886, 54.30428, 55.56258, 56.6066, 57.29723,
    58.68524, 58.74432, 57.17728, 55.50986, 52.687, 49.03281, 47.98659,
    46.7406, 44.42229, 43.40636, 45.28944, 47.52269, 48.2303, 46.90697,
    47.24905, 43.52259,
  55.74339, 58.87859, 59.45368, 54.66876, 59.17665, 66.35461, 68.37173,
    58.27041, 52.30606, 55.4288, 58.63389, 62.48159, 63.27113, 60.64411,
    58.21373, 55.89001, 50.57448, 45.22213, 44.21903, 43.07394, 41.25947,
    41.38415, 41.29479, 41.19946, 41.9221, 43.52176, 44.01402, 41.7571,
    39.06544, 37.03032,
  37.66483, 38.13866, 38.56223, 39.01054, 39.38291, 39.81248, 40.28693,
    40.81821, 41.36862, 42.06023, 43.47265, 43.66596, 42.0459, 42.55292,
    42.81182, 42.38265, 42.40035, 42.71311, 43.17072, 44.36252, 44.94094,
    44.30171, 44.95939, 46.13404, 46.67501, 46.13704, 48.89424, 48.71341,
    39.14342, 36.29435,
  43.26595, 44.08876, 44.20401, 45.2907, 45.57857, 45.93625, 46.70511,
    47.41257, 48.16085, 48.94333, 49.81948, 50.99284, 51.68683, 50.56787,
    50.06435, 50.35637, 49.34445, 49.38556, 49.90396, 50.38764, 49.9791,
    49.27957, 49.45665, 51.88737, 55.34587, 53.37795, 49.6809, 50.36972,
    40.05927, 37.25914,
  46.06913, 47.12919, 48.05375, 49.13527, 50.12827, 51.13077, 52.14834,
    53.29181, 54.48015, 55.52922, 56.46273, 57.51027, 58.40615, 59.75083,
    60.56585, 59.46984, 59.39132, 59.62839, 59.36071, 59.72402, 60.92289,
    62.07409, 62.07052, 62.38078, 63.40654, 60.83799, 55.58182, 49.66095,
    40.53621, 38.37612,
  51.37615, 53.02462, 54.59188, 56.27278, 57.92388, 59.73531, 60.77711,
    61.55468, 62.8813, 64.12003, 64.69431, 65.23929, 65.23985, 64.87018,
    66.77421, 67.76667, 65.44563, 62.87625, 63.05244, 63.52907, 65.62035,
    64.82471, 61.72434, 65.87051, 67.29057, 61.79684, 57.27866, 47.75951,
    40.13724, 36.73204,
  56.52156, 57.43243, 59.00266, 60.47602, 61.67811, 62.55864, 63.35586,
    64.39483, 66.19591, 67.54552, 67.56409, 67.81804, 67.74463, 68.1119,
    68.29634, 68.05391, 65.85725, 61.78912, 60.94255, 64.89985, 66.25842,
    59.36971, 59.22535, 61.45184, 63.93637, 61.83574, 55.50423, 55.07793,
    50.96749, 39.81879,
  63.1404, 65.94488, 68.43729, 70.91109, 71.29163, 71.24889, 72.55421,
    73.52465, 74.05756, 75.57452, 77.32927, 78.12089, 78.39535, 77.67744,
    77.28667, 77.92516, 78.49131, 76.44557, 65.61888, 64.57931, 60.79097,
    56.95139, 57.69211, 59.04427, 61.32854, 59.43345, 57.22586, 65.83535,
    59.23268, 38.5298,
  71.32516, 74.67617, 76.99894, 78.12285, 77.59325, 77.65538, 78.2667,
    78.31516, 77.75541, 77.20399, 75.25553, 71.46535, 66.86633, 66.41924,
    68.71021, 72.65536, 71.87967, 65.53349, 59.76472, 59.40668, 57.42661,
    56.2108, 56.91589, 59.41411, 59.296, 55.78965, 58.27273, 63.6183,
    53.98098, 36.331,
  72.31637, 74.62006, 76.03262, 77.07262, 75.714, 76.2658, 76.15921,
    69.51521, 65.37293, 65.13912, 64.27152, 63.39581, 62.78246, 63.62215,
    65.10956, 66.32871, 66.3318, 64.22379, 59.49161, 58.63913, 57.53699,
    57.58781, 59.50971, 60.84586, 57.83857, 56.09427, 62.23703, 60.77673,
    45.97893, 36.78888,
  77.80895, 79.66798, 80.85174, 80.85641, 79.9622, 80.52805, 77.72791,
    76.936, 78.95415, 80.37082, 81.16679, 81.58429, 81.85357, 83.04583,
    83.42001, 80.9977, 79.74643, 80.16409, 77.47178, 71.669, 68.21269,
    70.78079, 74.72065, 71.8811, 63.40704, 63.36757, 62.35764, 53.23713,
    40.00169, 36.40252,
  86.89039, 87.95073, 87.95203, 88.30454, 87.30962, 85.48179, 84.72513,
    85.56932, 85.86932, 86.51644, 86.97396, 87.641, 87.04738, 85.25079,
    83.31399, 82.99965, 82.06222, 80.60653, 76.51501, 72.56332, 71.67606,
    68.46654, 65.06284, 59.22131, 62.28468, 70.80727, 58.94764, 40.8598,
    36.38011, 34.84766,
  86.93177, 87.38209, 89.39549, 89.5376, 91.18143, 90.1096, 88.6461,
    87.65393, 87.06417, 87.50095, 87.2852, 81.95107, 81.11481, 78.80722,
    77.25289, 75.19215, 73.14905, 69.38667, 65.05773, 62.27708, 63.25974,
    58.4736, 50.17782, 46.43118, 47.45111, 46.5041, 40.48425, 36.10811,
    35.65811, 34.82048,
  88.54765, 84.87875, 87.88324, 89.38952, 88.82459, 87.46266, 86.51271,
    83.63902, 80.56649, 80.26973, 77.88211, 73.10402, 73.38806, 73.04767,
    69.19882, 65.97403, 61.93298, 59.15115, 56.42422, 55.42393, 56.54887,
    52.38367, 44.82848, 49.54556, 51.86359, 40.84472, 36.09241, 36.73014,
    36.20899, 35.32581,
  95.96207, 96.23927, 97.46004, 98.12633, 96.88731, 93.19606, 85.44109,
    82.08556, 82.88217, 80.00045, 80.65553, 79.89407, 80.00787, 80.21539,
    77.85785, 68.05318, 65.35126, 61.88958, 58.98215, 59.68739, 57.67305,
    49.8525, 45.54887, 45.87223, 46.30444, 39.43644, 36.78025, 36.96985,
    36.97318, 35.86261,
  88.7746, 89.08032, 89.03754, 87.24771, 86.00275, 85.45046, 85.66823,
    86.39463, 83.59906, 83.48341, 84.27191, 82.22141, 83.4015, 83.84689,
    81.33669, 78.9406, 76.19164, 74.07682, 72.06419, 66.81163, 56.01196,
    49.51633, 48.81752, 41.54722, 38.40694, 37.69091, 36.47019, 35.97717,
    36.15621, 35.64978,
  81.17397, 81.26916, 81.14764, 80.84488, 80.97961, 82.39842, 86.21232,
    87.6005, 84.76074, 84.5511, 83.9763, 83.39143, 83.15716, 81.95011,
    80.42262, 78.21124, 76.69241, 70.86649, 69.51999, 65.25277, 50.59139,
    47.22324, 41.03909, 38.85774, 37.71521, 37.31414, 36.46954, 35.84186,
    35.50229, 35.14587,
  82.70798, 83.36598, 83.83208, 83.72748, 83.60744, 84.69567, 85.77052,
    85.41974, 85.01169, 84.28589, 83.42585, 81.48592, 80.55493, 80.8111,
    79.17049, 74.74473, 69.72343, 61.85532, 58.10009, 54.12052, 43.16499,
    42.28235, 39.72754, 38.81535, 38.01133, 37.25054, 36.43447, 35.93381,
    35.52881, 35.10708,
  81.99832, 82.09563, 82.27432, 82.47007, 83.08597, 83.16634, 83.82166,
    84.61412, 84.13411, 83.527, 82.2445, 82.23165, 83.14111, 81.11873,
    75.91147, 69.38698, 63.30234, 57.46349, 57.27947, 54.65046, 42.09352,
    42.25869, 40.22256, 38.83148, 37.66161, 37.1677, 36.20633, 35.40281,
    35.21401, 35.02498,
  76.58813, 78.69449, 79.81699, 81.39666, 81.66252, 82.19306, 82.52759,
    83.05988, 83.5248, 82.68943, 82.74009, 83.01025, 81.96545, 80.82637,
    79.85579, 69.20598, 58.3124, 53.28933, 54.98101, 51.30165, 42.10504,
    41.27866, 39.58991, 38.49931, 36.81996, 36.28727, 35.94813, 35.09693,
    34.97711, 34.86437,
  75.96943, 75.30108, 74.09317, 74.89795, 77.13291, 78.42516, 80.02543,
    81.22709, 80.7598, 80.91575, 81.96085, 80.59494, 74.43163, 76.23492,
    76.41468, 73.81469, 72.32891, 70.5905, 70.03548, 63.66345, 51.02651,
    43.1832, 39.37629, 38.39474, 36.4725, 35.86105, 35.63046, 35.15324,
    34.95586, 34.84661,
  70.31618, 69.68181, 69.38695, 69.84762, 72.14577, 73.75936, 75.1828,
    76.31647, 77.458, 80.3221, 79.88891, 73.37838, 72.12334, 72.22709,
    71.29599, 68.87749, 67.9023, 66.77508, 64.92189, 62.33679, 55.36791,
    46.71792, 40.40346, 39.05888, 37.30748, 36.17798, 35.65316, 35.22008,
    34.95629, 34.85027,
  65.47483, 64.66798, 64.01894, 64.36337, 65.80167, 67.09634, 68.3271,
    69.48588, 70.97726, 72.61114, 69.39113, 64.53568, 65.1846, 64.23777,
    61.97429, 58.81185, 56.7952, 55.3775, 55.11763, 53.93523, 52.01051,
    49.85802, 45.18541, 41.29221, 38.54565, 36.79937, 35.71774, 35.26122,
    34.96851, 34.8699,
  64.84097, 61.39126, 60.3926, 60.22216, 60.97659, 60.95251, 61.83973,
    62.32315, 64.291, 64.28694, 59.36222, 56.67199, 57.02547, 55.98399,
    54.43632, 52.87553, 51.00836, 49.68882, 49.02622, 48.07487, 48.78365,
    49.65434, 48.04465, 46.77005, 42.20624, 37.93508, 35.92327, 35.53682,
    35.04494, 34.88348,
  63.71895, 61.64632, 59.6679, 59.26912, 60.85405, 61.41958, 60.60625,
    59.00915, 59.30114, 57.681, 53.71752, 53.91994, 54.18835, 53.85929,
    52.58021, 51.72003, 50.30995, 47.60952, 46.12652, 45.36295, 46.01311,
    46.77148, 44.7621, 44.99043, 44.47305, 40.21481, 36.87308, 36.44685,
    35.65642, 34.97419,
  70.51739, 68.66401, 68.15926, 68.35096, 68.61186, 68.17198, 68.6003,
    67.70771, 66.7599, 61.8245, 57.70749, 59.37829, 59.80279, 59.4814,
    57.71318, 55.51176, 53.37256, 50.5399, 47.37345, 46.01038, 46.05781,
    45.74226, 44.20634, 43.07122, 43.05746, 42.95792, 39.81308, 37.1458,
    36.35927, 35.33292,
  74.32257, 76.14244, 72.40208, 71.71293, 72.83239, 72.53915, 70.81989,
    69.57172, 69.80527, 66.14561, 61.2406, 62.66712, 62.85831, 61.52034,
    59.26049, 57.14093, 54.2354, 51.95267, 48.87534, 45.91717, 45.37607,
    44.79372, 43.44952, 42.31376, 41.29652, 42.18863, 42.21616, 39.48782,
    37.76563, 36.32222,
  81.70412, 85.43578, 83.12852, 79.6396, 77.89161, 76.50581, 76.54975,
    75.4865, 70.89245, 66.26347, 64.14601, 64.32929, 63.9767, 61.23362,
    57.79169, 55.63477, 53.56308, 51.62017, 49.34257, 46.81437, 46.34403,
    45.95374, 43.82412, 41.88374, 41.45415, 41.57031, 42.39433, 40.7659,
    37.37758, 36.0317,
  83.3757, 84.98833, 80.37831, 78.32759, 77.91339, 76.23167, 76.33141,
    73.97016, 68.31634, 65.22301, 64.90732, 64.76229, 63.72083, 61.22205,
    58.98656, 56.90247, 54.91726, 53.6466, 52.25121, 50.873, 51.80857,
    53.43377, 52.16902, 48.46053, 45.95807, 44.9815, 45.6633, 44.37324,
    38.13742, 35.04467,
  81.33985, 81.94864, 80.03353, 80.02947, 80.68359, 78.82635, 76.91978,
    72.75517, 67.51357, 67.48884, 67.512, 67.82359, 67.23314, 65.58836,
    64.37207, 62.28893, 59.8122, 58.47961, 57.67147, 57.09275, 56.82369,
    55.1631, 51.46037, 48.87369, 47.15171, 46.34325, 45.47207, 46.85751,
    44.1747, 36.90854,
  75.64364, 76.04596, 79.03737, 81.61777, 81.71223, 81.18362, 76.90586,
    70.00198, 67.35464, 68.17682, 67.81252, 67.73338, 67.69834, 67.80237,
    67.3727, 65.20773, 62.39493, 59.76231, 56.00483, 52.13269, 50.36682,
    48.29156, 45.79598, 44.08583, 43.71191, 43.47385, 42.59843, 41.00807,
    40.54931, 38.00024,
  74.89712, 76.3056, 77.0593, 76.74187, 77.04021, 79.029, 77.6101, 70.48724,
    66.96811, 68.85802, 69.92152, 70.24544, 69.08527, 67.29362, 64.44508,
    60.01472, 54.03001, 48.90813, 46.64942, 44.62021, 42.85044, 42.01667,
    41.20955, 40.46588, 40.08223, 40.09549, 39.54106, 38.02877, 36.42044,
    35.06699,
  32.75383, 32.83239, 32.89489, 32.96857, 32.99783, 33.05878, 33.14725,
    33.29459, 33.45905, 33.64804, 34.48772, 34.62218, 33.40466, 33.59368,
    33.74927, 33.41924, 33.41341, 33.6199, 33.88588, 34.65881, 35.13973,
    34.68333, 34.9347, 35.84612, 36.59701, 36.5267, 39.09105, 40.49104,
    35.19658, 33.429,
  34.33477, 34.52362, 34.31138, 34.678, 34.53116, 34.41683, 34.622, 34.81597,
    35.02374, 35.24113, 35.58177, 36.18751, 36.54185, 35.72097, 35.31944,
    35.56961, 35.15221, 35.51725, 36.28168, 37.05689, 37.33101, 37.34358,
    37.92015, 39.28799, 43.72837, 44.92966, 39.80679, 41.9825, 35.88532,
    34.08054,
  35.75648, 35.9217, 35.99146, 36.1377, 36.24732, 36.40544, 36.56487,
    36.78265, 37.04515, 37.25396, 37.51178, 38.0452, 38.43193, 39.01324,
    39.36572, 38.63558, 38.8648, 39.69576, 40.25867, 41.21325, 42.87215,
    44.78412, 45.7295, 45.27647, 49.19294, 51.4716, 43.1172, 41.35593,
    35.90617, 34.77095,
  38.96938, 39.38827, 39.86768, 40.4043, 40.948, 41.67654, 41.90762,
    41.79161, 42.05282, 42.46027, 42.73439, 43.28779, 43.40696, 42.98304,
    44.10052, 45.13076, 44.32616, 43.33161, 44.2083, 45.23075, 47.6114,
    48.44621, 46.45292, 51.10585, 53.38535, 46.41812, 45.33027, 40.0527,
    35.73338, 33.80501,
  43.78181, 43.86383, 44.45351, 45.06547, 45.46821, 45.64435, 45.77946,
    45.88157, 46.4907, 47.01106, 46.88801, 47.17774, 47.37013, 47.58165,
    47.68888, 47.79488, 46.74083, 45.25232, 45.32302, 49.95119, 51.90797,
    44.26834, 44.33419, 45.61669, 47.16716, 46.03796, 42.35588, 42.21779,
    41.56386, 35.7272,
  47.28657, 48.10898, 49.08462, 50.37303, 50.24868, 49.7589, 50.34403,
    50.72023, 50.76277, 51.42921, 52.4267, 54.78682, 57.08163, 56.17611,
    54.76135, 62.41435, 71.45371, 57.35936, 47.58468, 48.01626, 45.67598,
    42.54461, 43.28878, 44.43397, 46.48972, 45.1077, 47.80565, 63.01717,
    55.14782, 34.69121,
  51.59684, 53.06647, 54.49682, 56.09691, 56.61316, 57.04985, 58.51681,
    60.14608, 59.95724, 59.17779, 58.76213, 56.91085, 54.05175, 53.3201,
    56.76616, 61.95, 56.99347, 48.92303, 45.17444, 44.77229, 43.37651,
    42.60521, 43.29671, 45.53906, 46.26566, 42.59022, 51.45478, 67.90025,
    52.49652, 33.11381,
  56.29052, 57.93553, 59.35554, 60.69004, 60.27381, 61.29647, 62.10999,
    57.70351, 54.25737, 53.14299, 51.6574, 49.94238, 48.38673, 47.91901,
    47.90977, 47.95948, 47.32011, 45.97033, 43.28857, 42.87872, 42.17148,
    42.13977, 43.67378, 45.55831, 44.4282, 41.97688, 52.68714, 58.24548,
    39.62459, 33.77994,
  59.65858, 59.9615, 60.37959, 59.76907, 58.24091, 57.69689, 54.50401,
    52.26386, 52.00562, 51.62318, 50.89052, 50.08243, 49.7392, 52.81169,
    54.49866, 49.10021, 47.95265, 49.02492, 48.41715, 45.554, 43.61179,
    45.80316, 49.91136, 49.99472, 45.13248, 45.55174, 48.55363, 45.27169,
    35.87805, 33.61461,
  66.41292, 68.21035, 67.6263, 67.75416, 64.69915, 58.87558, 53.32347,
    54.60051, 55.2039, 56.86819, 58.83588, 61.90449, 61.59283, 58.10762,
    54.29963, 54.81921, 55.19862, 54.44493, 52.18423, 50.90938, 51.49002,
    50.83471, 49.83456, 45.94891, 53.19023, 66.56702, 52.64617, 36.63134,
    33.86627, 32.6203,
  79.80177, 79.29528, 79.13257, 78.22179, 77.79606, 75.41638, 70.83578,
    72.65125, 73.16745, 78.96878, 80.23071, 60.48179, 55.77998, 54.6651,
    53.93733, 53.70939, 53.8278, 52.87926, 51.19366, 50.16697, 51.7514,
    49.4699, 44.04119, 40.66898, 42.38364, 43.6475, 37.91575, 33.501,
    33.10836, 32.52695,
  86.68898, 82.04716, 85.45901, 85.95269, 85.07372, 83.37035, 82.09314,
    78.65096, 69.75459, 69.19911, 65.3776, 57.49526, 58.55814, 57.72897,
    53.13608, 52.27723, 49.99733, 48.6897, 47.05625, 46.28707, 47.5222,
    45.14274, 39.03822, 42.97438, 45.4653, 36.04817, 33.20729, 33.58653,
    33.38424, 32.80948,
  94.74696, 94.79787, 97.33439, 96.61028, 94.40181, 89.50245, 80.67873,
    75.48769, 75.90202, 70.42738, 69.63829, 63.86414, 64.56548, 64.25024,
    55.51169, 50.47198, 48.48778, 46.88519, 45.30178, 46.33535, 46.32653,
    41.95925, 38.41278, 41.27503, 42.95209, 35.02383, 33.63066, 33.74694,
    33.83072, 33.14534,
  92.1656, 94.70402, 92.6151, 88.81004, 85.08827, 82.41626, 81.10993,
    80.7879, 78.12846, 76.8958, 78.07116, 76.6242, 77.54475, 77.85318,
    76.41611, 58.93074, 49.48127, 50.26207, 50.49509, 49.41869, 44.3511,
    42.94437, 45.39531, 38.02676, 35.20015, 34.34941, 33.59571, 33.24001,
    33.38656, 33.02195,
  82.51662, 81.4593, 79.72799, 77.78448, 76.31508, 77.90297, 83.28607,
    82.86137, 79.39684, 78.49302, 77.18613, 75.56596, 68.04364, 70.92904,
    70.9054, 55.28559, 53.25618, 50.78247, 51.39559, 52.33485, 47.92899,
    41.89981, 36.77258, 34.9365, 34.25619, 34.29351, 33.63338, 33.14494,
    32.96289, 32.73286,
  78.26775, 77.76443, 77.52702, 76.822, 76.26027, 76.82561, 77.45057,
    76.8501, 75.93088, 72.2738, 68.96163, 63.62837, 59.80229, 59.97133,
    55.79511, 51.87588, 50.2663, 46.53838, 45.44173, 44.14189, 38.0584,
    36.58607, 34.81833, 34.47275, 34.42067, 34.15531, 33.64429, 33.20678,
    32.93156, 32.68733,
  76.98265, 75.49762, 74.25047, 73.29457, 72.68594, 71.35789, 70.32724,
    69.39625, 67.27232, 65.21219, 60.75948, 60.32987, 62.23322, 56.71043,
    51.74846, 48.58455, 45.79735, 42.98199, 43.92014, 43.04301, 35.80238,
    36.09649, 35.24612, 34.52775, 34.16837, 34.12843, 33.51407, 32.92488,
    32.7808, 32.6539,
  68.16875, 67.7499, 65.98274, 65.02822, 63.68736, 63.08821, 62.46244,
    62.06227, 61.72078, 59.1383, 59.22644, 60.49981, 57.57408, 54.71922,
    53.42117, 48.01695, 42.46245, 40.00859, 42.27362, 41.21403, 35.83795,
    35.90197, 35.27242, 34.70832, 33.80404, 33.60026, 33.33936, 32.74335,
    32.63809, 32.55802,
  65.72453, 64.13266, 60.77435, 58.54093, 57.76596, 56.79223, 56.28267,
    56.06711, 54.97097, 54.04582, 55.0453, 53.03954, 47.87754, 47.66941,
    47.17023, 45.64871, 45.77735, 46.63591, 48.84468, 47.87455, 41.90928,
    37.502, 35.17844, 34.80057, 33.63271, 33.25127, 33.10261, 32.75313,
    32.61237, 32.54065,
  61.74171, 59.61731, 56.60133, 54.018, 53.21271, 52.45506, 51.85091,
    51.3117, 50.89709, 52.37963, 52.25484, 47.77813, 46.47223, 46.37249,
    45.89111, 45.07676, 45.95023, 47.21428, 47.94247, 47.81121, 44.48118,
    39.40898, 35.42363, 34.93095, 34.03343, 33.39851, 33.08805, 32.78721,
    32.60799, 32.53942,
  58.22422, 56.23292, 53.34485, 51.13727, 50.18439, 49.59693, 49.21239,
    48.99127, 49.48216, 51.0214, 49.47967, 46.47193, 47.30424, 47.03246,
    45.68599, 43.88499, 43.05702, 42.50065, 42.44564, 41.79546, 40.55069,
    39.56119, 37.65068, 35.97538, 34.65766, 33.75613, 33.13464, 32.80589,
    32.61781, 32.55315,
  57.89867, 54.82819, 52.34701, 50.58796, 49.80243, 48.86104, 48.68703,
    48.50889, 49.86174, 50.47697, 47.49875, 45.45174, 45.48542, 44.34907,
    42.67067, 41.19656, 39.84013, 38.95354, 38.58114, 37.93711, 39.02139,
    39.9735, 38.42731, 38.80864, 36.6727, 34.33912, 33.20357, 32.95696,
    32.65838, 32.55845,
  56.92419, 55.12169, 52.42377, 50.88385, 51.10357, 50.98421, 50.04126,
    48.57482, 48.69021, 47.4568, 44.06643, 43.23073, 42.68255, 41.72739,
    40.28093, 39.62795, 39.02106, 37.68415, 37.12537, 36.77378, 37.88566,
    38.68658, 36.59031, 37.58564, 37.77019, 35.51797, 33.63885, 33.49557,
    33.04947, 32.61397,
  57.10436, 55.77008, 54.34998, 53.56829, 52.94802, 51.80423, 51.32284,
    50.48217, 49.988, 46.59907, 42.8452, 42.91097, 42.73747, 42.37346,
    41.3911, 40.50163, 40.0396, 38.952, 37.43624, 36.83799, 36.92036,
    36.83257, 36.15028, 35.98254, 36.55638, 36.91856, 35.36569, 33.93087,
    33.47309, 32.82173,
  56.43777, 56.60229, 53.63243, 52.15306, 51.939, 51.06113, 49.66321,
    48.90901, 49.41741, 46.79329, 42.9305, 43.37908, 43.53922, 42.99671,
    42.03809, 41.3673, 40.40156, 39.76318, 38.50989, 37.0726, 36.92582,
    36.88864, 36.4644, 35.8099, 35.2905, 36.31423, 36.5776, 35.0723,
    34.25151, 33.36506,
  57.25549, 58.41181, 56.61547, 53.94675, 51.8833, 50.55571, 50.80562,
    51.12181, 49.12351, 46.04215, 44.43565, 44.70016, 44.80268, 43.46212,
    41.60651, 40.80563, 40.18572, 39.69736, 38.82672, 37.38079, 37.24184,
    37.28027, 36.25957, 35.40285, 35.37966, 35.77233, 36.7054, 35.89755,
    34.05248, 33.19878,
  58.42051, 58.56519, 55.16054, 52.85881, 51.66594, 50.23452, 50.8569,
    50.56277, 47.54525, 45.31925, 45.12799, 45.05303, 44.36584, 42.83941,
    41.4401, 40.38031, 39.55121, 39.24654, 38.6191, 37.58937, 38.15553,
    39.70011, 39.9785, 38.5512, 37.5145, 37.36266, 38.41894, 38.04247,
    34.4168, 32.5941,
  57.79188, 56.76449, 54.39071, 53.50368, 53.16098, 51.7712, 51.22514,
    49.24374, 45.65953, 44.96181, 44.56311, 44.26515, 43.52261, 42.33576,
    41.74826, 40.99144, 40.07503, 40.03576, 40.34164, 40.59811, 41.34658,
    41.47942, 40.13047, 38.892, 38.18017, 38.0607, 37.91251, 39.22488,
    37.82488, 33.70002,
  55.43647, 54.02747, 54.23833, 54.74252, 54.39417, 54.22563, 51.77181,
    47.09679, 44.61871, 44.38779, 43.44889, 42.90279, 42.64133, 42.7406,
    43.28828, 43.44713, 43.29839, 43.33846, 42.22321, 40.54222, 40.08451,
    39.23385, 37.88203, 37.04379, 36.98752, 37.08183, 36.82275, 36.24302,
    36.3028, 34.46867,
  54.80283, 54.62057, 54.17431, 53.01103, 52.36406, 53.70421, 53.46759,
    48.60761, 45.65391, 46.34768, 46.85368, 47.26123, 47.0218, 46.48556,
    45.92088, 44.98204, 42.84439, 40.60435, 39.53329, 38.24658, 37.16865,
    36.66032, 36.20313, 35.81191, 35.5788, 35.68378, 35.43983, 34.61,
    33.7456, 32.80387,
  28.8234, 28.8584, 28.89778, 28.94344, 28.93984, 28.94597, 28.9897,
    29.03547, 29.14497, 29.2823, 30.01303, 30.12748, 29.14259, 29.28786,
    29.39394, 29.0976, 29.03301, 29.10459, 29.18554, 29.67538, 29.93793,
    29.45977, 29.46478, 30.06391, 30.53399, 30.4165, 32.69688, 34.07367,
    30.59042, 29.40069,
  29.38405, 29.46318, 29.25124, 29.52097, 29.41633, 29.27474, 29.35969,
    29.47126, 29.61155, 29.77442, 30.07864, 30.57587, 30.83912, 30.17585,
    29.83944, 29.93547, 29.51036, 29.63779, 30.08757, 30.55841, 30.60201,
    30.3263, 30.65831, 31.51734, 35.55276, 36.8976, 33.20343, 35.36616,
    31.12945, 29.81423,
  29.51727, 29.54925, 29.5544, 29.59119, 29.59145, 29.62414, 29.65928,
    29.76098, 29.89533, 29.98736, 30.11263, 30.46866, 30.70727, 31.13234,
    31.32704, 30.67361, 30.72175, 31.23809, 31.53867, 32.07264, 33.21801,
    34.62624, 35.75897, 35.45503, 40.00047, 42.92678, 35.53828, 35.16077,
    31.23545, 30.36317,
  30.17429, 30.28084, 30.5156, 30.77477, 31.09464, 31.56157, 31.65295,
    31.50455, 31.60346, 31.85067, 31.90594, 32.20853, 32.22951, 31.88781,
    32.88726, 33.95784, 33.54816, 32.91893, 33.64248, 34.50708, 36.757,
    37.98748, 36.74196, 41.69783, 44.2058, 38.223, 37.62846, 34.20904,
    31.11186, 29.74296,
  31.98381, 31.92791, 32.31082, 32.76513, 33.06503, 33.20469, 33.31567,
    33.32225, 33.77361, 34.04809, 33.76321, 33.80619, 33.92508, 34.29768,
    34.93408, 35.57796, 35.16186, 34.83667, 35.31484, 40.10382, 42.11913,
    35.87807, 35.87292, 37.31384, 38.72139, 37.4323, 34.96744, 34.79141,
    34.93262, 31.17842,
  33.7745, 34.24141, 35.03871, 35.97477, 35.79843, 35.38012, 35.75191,
    35.90144, 35.80404, 36.16082, 36.63517, 38.38922, 40.31036, 40.29521,
    39.37313, 47.12508, 56.65916, 45.97299, 38.05975, 39.23035, 37.55553,
    34.58469, 34.97744, 35.61598, 37.48756, 36.39848, 39.34674, 53.16133,
    47.05179, 30.34378,
  36.01047, 36.82124, 37.85555, 38.94611, 39.2366, 39.60366, 41.04334,
    42.94387, 43.42926, 43.35205, 43.66132, 42.83155, 41.17775, 40.68452,
    45.44651, 52.61525, 48.36891, 40.0852, 37.01985, 36.45621, 35.15901,
    34.48372, 34.94489, 36.76872, 37.75283, 34.62741, 43.86341, 60.18934,
    45.94922, 29.22773,
  39.073, 40.38691, 41.90377, 43.47011, 43.8165, 45.64692, 47.7529, 45.73948,
    43.77633, 43.41195, 42.4921, 40.93629, 39.29361, 38.59922, 39.20813,
    39.86427, 38.71318, 37.338, 35.4283, 35.01735, 34.42595, 34.23452,
    35.38869, 36.95474, 36.41598, 34.09452, 45.99235, 52.2029, 34.63023,
    30.04948,
  44.36761, 45.47714, 46.66449, 47.05613, 46.86149, 47.40279, 45.69439,
    44.04851, 43.66401, 43.03549, 41.84715, 40.36082, 39.2007, 41.29296,
    42.3853, 38.34445, 37.81847, 38.96297, 38.59891, 36.35591, 34.70583,
    36.11855, 39.54865, 39.72837, 36.17583, 36.54022, 40.92438, 39.60749,
    32.10345, 29.98724,
  50.11879, 52.28188, 52.66669, 53.07773, 51.53849, 47.29861, 42.76118,
    42.86222, 42.63026, 42.85176, 43.89796, 46.54194, 46.46284, 43.91654,
    40.97137, 41.04073, 41.64791, 41.37501, 39.97571, 39.56348, 40.08981,
    40.29727, 40.45025, 37.99524, 44.69352, 55.64271, 45.039, 32.69481,
    30.37008, 29.01426,
  72.13411, 73.76826, 66.84904, 58.51235, 56.00089, 52.32257, 48.37848,
    50.75967, 52.07763, 60.83151, 67.52924, 46.885, 41.51297, 40.20359,
    39.31072, 39.84585, 41.40196, 40.95982, 39.70637, 39.50444, 42.03057,
    41.09116, 37.1025, 34.46199, 37.65702, 40.44464, 34.55304, 29.89537,
    29.38437, 28.88032,
  81.43624, 76.47314, 79.43188, 81.11827, 81.10856, 68.42857, 68.17508,
    61.3924, 50.91559, 54.06509, 53.01278, 41.22498, 42.263, 42.31236,
    39.03566, 39.89328, 38.99257, 38.56243, 37.63299, 37.66634, 40.2667,
    38.73409, 33.51902, 37.08775, 39.01411, 31.81977, 29.33852, 29.74848,
    29.61645, 29.07375,
  84.98205, 85.13738, 90.28935, 92.32464, 93.11361, 90.02009, 76.75417,
    53.36385, 53.51467, 49.30974, 47.70189, 42.74122, 45.41693, 46.17023,
    40.3968, 39.53703, 38.87101, 37.82664, 36.79015, 38.58265, 39.72443,
    36.0836, 32.87346, 37.02507, 38.41365, 30.91471, 29.65015, 29.86931,
    30.04776, 29.37283,
  87.51759, 92.96595, 92.62613, 90.81681, 87.99435, 84.10661, 80.24912,
    79.95334, 71.56354, 67.83638, 76.43176, 71.08972, 71.26089, 68.1302,
    58.41066, 46.04251, 39.06995, 40.36192, 41.43055, 41.88425, 38.34311,
    37.15379, 39.05154, 34.03087, 31.49723, 30.26238, 29.65268, 29.41421,
    29.69179, 29.29837,
  79.93634, 79.76942, 74.09169, 69.47739, 64.6414, 75.50893, 82.73075,
    83.16412, 80.6861, 80.23485, 76.94832, 60.94075, 49.38625, 54.10705,
    57.42207, 43.15131, 42.94281, 42.18422, 45.23759, 46.69305, 41.37598,
    36.92365, 32.99867, 30.80248, 30.04136, 30.36432, 29.7605, 29.32877,
    29.26363, 29.04613,
  63.21405, 60.76721, 59.34966, 58.09665, 58.50467, 63.05431, 67.34575,
    64.26332, 60.83472, 57.32415, 52.72692, 46.40601, 43.35591, 45.61242,
    44.47478, 42.12432, 42.90911, 40.63411, 41.22877, 40.68787, 34.40374,
    32.05898, 30.22767, 30.06596, 30.33933, 30.28196, 29.85685, 29.43999,
    29.21839, 28.99078,
  58.10044, 56.31847, 55.32707, 55.04136, 55.2832, 54.51722, 53.46214,
    52.6964, 50.83871, 48.47791, 44.72349, 45.27191, 48.693, 45.21434,
    41.96008, 40.99782, 39.85059, 37.59664, 39.53254, 38.57156, 31.09457,
    31.30074, 30.77333, 30.22533, 30.1394, 30.27246, 29.75484, 29.21075,
    29.1054, 28.96388,
  53.94886, 53.43932, 52.20316, 51.55282, 50.38668, 49.55701, 48.92556,
    48.47069, 47.58668, 45.59977, 45.61563, 47.90556, 46.36324, 44.54627,
    45.02613, 41.57914, 36.89973, 34.53751, 37.73869, 36.89177, 31.37481,
    31.56217, 31.1474, 30.61762, 29.84892, 29.86884, 29.57835, 29.04314,
    28.9644, 28.88953,
  53.14991, 51.97163, 49.28307, 47.36539, 46.55778, 45.68896, 45.32264,
    45.28661, 44.37963, 43.62195, 45.23166, 43.86965, 38.70751, 38.5744,
    38.66812, 37.40667, 37.40622, 38.26937, 41.5387, 41.11454, 35.54657,
    32.65841, 31.38346, 30.84747, 29.79989, 29.53061, 29.3918, 29.05397,
    28.92262, 28.86943,
  50.83631, 49.15084, 46.6509, 44.63839, 44.13836, 43.68705, 43.31627,
    42.9217, 42.40112, 43.77103, 43.43581, 38.31792, 35.6466, 35.39033,
    35.17429, 34.58823, 36.04056, 38.10922, 40.32342, 41.45189, 38.61509,
    34.61055, 31.7137, 31.00964, 30.19097, 29.62216, 29.36113, 29.07403,
    28.91715, 28.87199,
  47.95564, 46.88482, 45.00896, 43.12836, 42.45023, 42.00961, 41.49458,
    40.84674, 40.77659, 41.91959, 39.41514, 35.08356, 35.14223, 35.41325,
    35.12622, 34.37678, 34.54546, 34.91182, 36.03661, 36.44538, 35.76418,
    35.23412, 33.72843, 31.91398, 30.64876, 29.8891, 29.37873, 29.08625,
    28.94435, 28.8805,
  47.02336, 45.69691, 43.55406, 42.07597, 41.25918, 40.17131, 39.64604,
    39.09317, 40.20181, 40.50513, 36.92783, 34.51126, 34.86507, 34.78706,
    34.42028, 34.01388, 33.40422, 33.0101, 33.03253, 32.67751, 33.86852,
    34.75121, 34.41075, 34.84877, 32.78924, 30.50854, 29.46365, 29.24087,
    28.97874, 28.89166,
  46.03163, 44.49375, 41.95591, 40.45574, 40.66352, 40.74829, 40.17353,
    39.27491, 40.22148, 39.21332, 35.55424, 34.47357, 34.29465, 34.06448,
    33.49302, 33.58419, 33.33221, 32.2201, 31.71287, 31.49866, 32.84103,
    33.42283, 32.28261, 33.80485, 34.08297, 31.66977, 29.81432, 29.70639,
    29.3149, 28.93463,
  44.90879, 43.32514, 42.15402, 41.75763, 41.68926, 41.45722, 41.93806,
    42.28616, 43.04998, 39.76677, 35.37035, 34.90385, 34.67017, 34.72343,
    34.41043, 34.15951, 34.26255, 33.41865, 31.99843, 31.66031, 32.07664,
    32.06947, 31.5694, 31.74791, 32.862, 33.17881, 31.41529, 30.06684,
    29.69043, 29.11283,
  44.25745, 44.65079, 42.17093, 41.37466, 41.86757, 41.84348, 41.35004,
    41.52721, 42.96591, 39.91977, 35.21239, 34.87131, 34.93052, 34.8752,
    34.69165, 34.75244, 34.44647, 34.21141, 33.01908, 31.63603, 31.83329,
    32.07297, 31.87256, 31.24394, 30.83774, 32.09133, 32.28629, 30.93007,
    30.46584, 29.55899,
  45.25026, 46.82084, 45.54335, 43.63855, 42.20614, 41.23521, 42.14909,
    43.23038, 41.76579, 38.38274, 35.77532, 35.50094, 35.75154, 35.07523,
    34.20404, 34.20421, 34.06895, 34.0271, 33.29307, 31.91102, 32.21227,
    32.51531, 31.49799, 30.73434, 30.63244, 31.11332, 32.39254, 31.6964,
    30.28583, 29.39564,
  46.74863, 47.70752, 44.65921, 42.61492, 41.58926, 40.52612, 41.84148,
    42.47955, 39.6558, 36.96958, 36.11944, 35.84275, 35.53684, 34.67993,
    34.13342, 33.88149, 33.59398, 33.67114, 33.03397, 31.81264, 32.53789,
    34.29985, 34.70713, 33.30142, 32.33242, 32.36101, 33.90285, 33.71738,
    30.46234, 28.85483,
  46.22871, 45.71439, 43.53898, 42.81712, 42.82159, 41.97103, 42.35304,
    41.09132, 37.69808, 36.69207, 35.89471, 35.46422, 34.99873, 34.34708,
    34.3789, 34.10033, 33.47654, 33.51608, 33.64218, 33.58508, 35.07685,
    35.90586, 34.93509, 33.54004, 32.72904, 32.83209, 33.0318, 34.85772,
    33.47182, 29.76494,
  43.41566, 42.24697, 42.69777, 43.82286, 44.38728, 45.16911, 43.60357,
    39.6063, 37.23442, 36.70828, 35.11032, 33.83717, 33.20621, 33.47947,
    34.49369, 35.03761, 35.24473, 35.84698, 34.98734, 33.59158, 33.76899,
    33.38098, 32.23419, 31.49751, 31.5696, 31.97266, 32.00087, 31.86931,
    32.42641, 30.45778,
  42.35987, 42.48938, 42.64503, 42.20913, 42.19796, 44.5416, 44.8732,
    40.04478, 37.05793, 37.11106, 36.74398, 36.30233, 35.95187, 36.26428,
    36.81414, 36.78928, 35.60675, 34.23254, 33.39513, 32.21027, 31.48483,
    31.19094, 30.91915, 30.69992, 30.69421, 31.1189, 31.11563, 30.4905,
    29.95451, 29.14831,
  25.62791, 25.65708, 25.69319, 25.73092, 25.72091, 25.71124, 25.72384,
    25.76323, 25.84065, 25.95178, 26.80931, 26.95063, 25.90379, 26.05731,
    26.17785, 25.84199, 25.75684, 25.80329, 25.83739, 26.34599, 26.60337,
    26.08632, 26.05385, 26.60944, 26.93465, 26.63447, 29.06579, 30.86232,
    27.60512, 26.35373,
  26.02328, 26.09645, 25.87528, 26.13947, 25.98792, 25.83521, 25.9102,
    25.9936, 26.11244, 26.27325, 26.64142, 27.18401, 27.46835, 26.79659,
    26.41842, 26.47836, 25.98477, 26.04055, 26.45141, 26.91814, 26.89699,
    26.44556, 26.49742, 27.34804, 31.01506, 31.87787, 29.52434, 32.53886,
    28.22113, 26.83483,
  25.97468, 26.00287, 25.98486, 26.02746, 25.9727, 25.95601, 25.99751,
    26.0845, 26.19545, 26.26194, 26.35516, 26.76226, 27.04548, 27.47083,
    27.58973, 26.74999, 26.6763, 27.05061, 27.10981, 27.41714, 28.31384,
    29.60795, 30.60012, 30.41648, 34.93573, 37.75602, 31.93892, 32.34499,
    28.22586, 27.41208,
  26.0844, 26.11705, 26.30016, 26.47202, 26.74637, 27.23291, 27.3118,
    27.09285, 27.15224, 27.41285, 27.47772, 27.7946, 27.68494, 27.22927,
    28.21114, 29.19475, 28.6004, 27.64605, 27.97819, 28.51567, 30.96766,
    32.42626, 31.39431, 36.16013, 38.45128, 34.25179, 34.75849, 31.7226,
    28.18584, 26.71836,
  26.84974, 26.5982, 26.87177, 27.22316, 27.55096, 27.75147, 27.77563,
    27.68223, 28.19196, 28.54728, 28.22269, 28.15641, 28.10737, 28.39436,
    29.1481, 29.76484, 29.08682, 28.44736, 29.03193, 33.36078, 35.31449,
    30.54059, 30.46233, 32.39595, 34.22633, 33.48865, 31.61385, 31.672,
    32.31026, 28.37876,
  27.30601, 27.47228, 28.19817, 29.14364, 29.01487, 28.56996, 28.73901,
    28.62443, 28.2799, 28.37153, 28.52631, 30.31103, 32.54572, 32.55597,
    32.04193, 39.10721, 47.06996, 38.37952, 32.13354, 33.89047, 32.37271,
    29.19013, 29.61813, 30.46221, 32.85125, 32.33998, 33.9597, 45.9227,
    42.60459, 27.78111,
  28.18088, 28.57402, 29.348, 30.22143, 30.31474, 30.29082, 31.25136,
    32.93097, 33.34114, 33.21677, 33.78857, 33.51991, 32.36665, 32.49602,
    37.30522, 44.69192, 42.34224, 34.5784, 31.7114, 31.39853, 29.96551,
    29.03623, 29.53039, 31.81118, 33.25974, 30.68295, 39.06361, 54.48293,
    43.12482, 26.42428,
  29.31026, 29.9026, 30.98579, 32.20969, 32.3726, 34.53077, 37.06938,
    35.11578, 33.45155, 33.49369, 33.16099, 32.08839, 30.972, 31.11095,
    32.8889, 34.43897, 33.38309, 31.97266, 30.17077, 29.82841, 29.18012,
    28.90286, 30.20698, 32.52588, 32.19026, 30.31559, 42.08809, 48.33367,
    32.49467, 26.67425,
  32.31735, 32.92028, 34.24034, 34.84753, 35.271, 37.04681, 36.12538,
    34.53321, 34.38461, 34.15165, 33.16892, 31.86048, 31.06238, 34.13652,
    36.33334, 32.60486, 32.12889, 33.678, 33.58542, 31.25931, 29.20488,
    30.59101, 34.66756, 35.56475, 31.82043, 32.22869, 38.4304, 37.18344,
    28.49692, 26.68654,
  36.85897, 39.14123, 40.98662, 42.82428, 42.19625, 38.4718, 34.13894,
    34.02866, 33.49995, 33.11592, 34.03458, 37.42963, 38.53623, 37.20142,
    34.95957, 34.97158, 35.82859, 36.32244, 34.73701, 32.94717, 33.14025,
    33.65028, 34.48668, 32.63429, 38.00209, 48.52354, 40.95781, 29.53375,
    27.06987, 25.88753,
  52.11366, 54.53913, 50.32208, 45.10394, 43.08984, 41.41758, 37.46353,
    39.48418, 41.222, 48.63993, 53.61486, 38.4549, 33.97694, 33.14944,
    32.49313, 33.25804, 34.4614, 34.40887, 33.17717, 32.8173, 35.49291,
    35.11004, 31.9006, 29.69488, 33.48269, 37.35408, 31.6711, 26.58848,
    26.22729, 25.7351,
  68.83602, 55.27574, 57.59452, 58.8816, 57.95432, 50.42302, 52.70378,
    49.33401, 41.35835, 45.25586, 44.99763, 32.60813, 33.36034, 34.16831,
    32.23611, 32.71932, 32.14214, 32.03818, 31.58147, 31.94325, 34.89362,
    33.81482, 29.33519, 32.61112, 34.53746, 28.43042, 26.13192, 26.50644,
    26.39729, 25.90017,
  78.64268, 74.82102, 90.48232, 93.34669, 95.88964, 86.68104, 64.92475,
    43.59138, 42.76912, 39.87991, 37.22855, 31.93218, 35.75356, 37.87223,
    33.66581, 32.749, 32.85834, 32.075, 31.25901, 33.32517, 34.9164,
    31.72572, 28.87886, 33.36902, 34.76024, 27.59445, 26.34014, 26.63866,
    26.862, 26.18351,
  84.16695, 94.96472, 96.53934, 96.16403, 85.47375, 74.23282, 68.46291,
    62.43415, 53.31253, 48.59109, 56.61462, 54.75308, 56.57523, 54.95422,
    48.83979, 39.36385, 33.42469, 34.77139, 35.9294, 37.02411, 34.10012,
    32.72419, 34.5309, 30.80404, 28.4526, 26.91137, 26.39224, 26.22861,
    26.55561, 26.13894,
  63.47718, 68.94428, 64.66087, 60.13338, 53.34032, 59.08934, 79.35889,
    75.49248, 67.07287, 67.43517, 64.3382, 51.8972, 42.24619, 47.10704,
    49.25801, 36.7737, 36.88755, 36.93983, 40.35761, 41.61172, 36.44473,
    33.08113, 30.13784, 27.65209, 26.70877, 27.04955, 26.49345, 26.13986,
    26.12086, 25.8968,
  50.31807, 48.46804, 46.64185, 44.46373, 44.15396, 49.32536, 55.57879,
    53.36886, 50.64845, 48.95958, 45.76205, 39.03831, 34.85657, 38.40178,
    38.40155, 36.0425, 37.70043, 36.1935, 37.61293, 37.39097, 31.32237,
    28.82095, 26.90808, 26.76941, 27.10313, 27.02861, 26.58994, 26.2382,
    26.07154, 25.82586,
  45.20789, 42.75277, 41.33601, 41.01293, 42.09298, 42.96175, 43.15425,
    43.08441, 41.87665, 40.06314, 36.23127, 36.09711, 40.28526, 38.26937,
    36.1525, 36.05151, 35.71415, 33.85225, 35.71802, 34.68568, 27.83065,
    27.80757, 27.40492, 26.91971, 26.8698, 27.00571, 26.52971, 26.02931,
    25.9728, 25.81928,
  40.45921, 39.80333, 39.35582, 39.88773, 39.99601, 40.22087, 40.06722,
    39.70295, 39.00502, 36.32465, 36.12532, 39.34114, 39.50606, 38.56498,
    39.67252, 37.36121, 33.23858, 30.93557, 33.96436, 33.04447, 27.85542,
    28.12904, 27.79961, 27.25862, 26.57855, 26.65348, 26.37016, 25.87621,
    25.82759, 25.75248,
  40.77023, 40.81753, 39.36871, 38.44092, 38.18501, 37.61192, 37.21421,
    36.81695, 35.69904, 34.72306, 37.1011, 37.40083, 33.4319, 33.969,
    34.73866, 33.58302, 33.15544, 33.69203, 36.73797, 36.16066, 31.21111,
    29.10693, 28.10245, 27.55248, 26.59105, 26.35949, 26.19789, 25.88056,
    25.79238, 25.7266,
  41.29771, 40.80548, 38.85823, 36.94036, 36.48648, 36.01247, 35.59803,
    35.12427, 34.65453, 36.45121, 37.23065, 33.12221, 30.77255, 30.92942,
    30.8056, 30.09285, 31.37902, 33.46668, 35.88743, 37.0048, 34.47987,
    30.98565, 28.44676, 27.77748, 26.98224, 26.43979, 26.15859, 25.89781,
    25.78794, 25.72561,
  40.35852, 39.62408, 37.61876, 35.91524, 35.34534, 35.14305, 34.89106,
    34.4673, 34.60034, 36.11628, 34.06264, 29.82104, 30.01345, 30.46223,
    30.23163, 29.48219, 29.78509, 30.5248, 32.01418, 32.74683, 32.27894,
    31.6844, 30.20908, 28.4937, 27.39241, 26.68919, 26.17805, 25.92053,
    25.81258, 25.73462,
  40.37673, 38.55422, 36.82188, 35.61841, 35.15871, 34.52349, 34.24037,
    33.69002, 34.5358, 34.6138, 30.96705, 28.66893, 29.42006, 29.76057,
    29.64054, 29.42705, 29.12277, 29.02332, 29.27659, 29.09411, 30.18064,
    31.02192, 31.02694, 31.35585, 29.45555, 27.28741, 26.31283, 26.0716,
    25.85912, 25.75301,
  39.51535, 38.18616, 36.2046, 35.00339, 35.27525, 35.39204, 34.76009,
    33.4899, 33.98273, 32.75264, 29.18311, 28.52971, 29.00784, 29.26018,
    29.06643, 29.45311, 29.33997, 28.37528, 27.97485, 27.89248, 29.2414,
    29.71509, 29.04868, 30.64898, 30.77935, 28.29394, 26.59278, 26.49093,
    26.13823, 25.79094,
  38.84872, 37.6601, 36.51015, 35.99268, 35.85549, 35.59349, 35.72206,
    35.47142, 35.87957, 32.81438, 28.98376, 29.21768, 29.74401, 30.22827,
    30.17019, 30.19815, 30.29718, 29.42476, 28.27124, 28.12699, 28.57216,
    28.52819, 28.17214, 28.57281, 29.7233, 29.81818, 28.06787, 26.81236,
    26.48011, 25.93103,
  38.05425, 38.31021, 36.10089, 35.11698, 35.41019, 35.3367, 34.86429,
    34.89581, 36.20458, 33.27069, 29.17605, 29.5479, 30.24226, 30.6254,
    30.65898, 30.75508, 30.54196, 30.31553, 29.14674, 27.95316, 28.2738,
    28.54852, 28.394, 27.7865, 27.51239, 28.76507, 28.84967, 27.54824,
    27.22438, 26.332,
  38.13932, 39.61564, 38.34733, 36.60785, 35.38831, 34.55911, 35.43044,
    36.44714, 35.34595, 32.12806, 29.83491, 30.23767, 31.05948, 30.76003,
    30.14329, 30.29676, 30.1947, 30.13977, 29.39491, 28.16229, 28.61521,
    28.9336, 27.97837, 27.2291, 27.10131, 27.70367, 29.02637, 28.26716,
    27.10069, 26.20739,
  38.91779, 40.25052, 37.57955, 35.69724, 34.90105, 34.10366, 35.50274,
    36.23146, 33.49074, 30.73895, 30.15205, 30.50811, 30.80828, 30.36067,
    30.02916, 29.91752, 29.71032, 29.8031, 29.15371, 28.03313, 28.85829,
    30.44255, 30.60009, 29.27257, 28.57941, 28.76608, 30.50602, 30.26664,
    27.19521, 25.69836,
  38.41343, 38.36946, 36.41862, 35.77349, 36.11158, 35.63236, 36.33873,
    35.03733, 31.45328, 30.30024, 29.91795, 30.18887, 30.34562, 30.11688,
    30.37899, 30.20554, 29.59738, 29.54626, 29.57254, 29.46378, 30.96772,
    31.77227, 30.86968, 29.5564, 29.04198, 29.24228, 29.65385, 31.50003,
    29.94177, 26.45742,
  35.9056, 34.92971, 35.42452, 36.63924, 37.65089, 38.8834, 37.65538,
    33.60466, 30.90712, 30.3289, 29.24789, 28.69945, 28.67995, 29.25581,
    30.33604, 30.9438, 31.16199, 31.50102, 30.55882, 29.38669, 29.69817,
    29.41306, 28.36343, 27.77271, 27.99026, 28.43595, 28.5441, 28.64983,
    29.2591, 27.14045,
  35.07014, 35.20491, 35.5492, 35.47673, 35.88139, 38.52819, 38.96181,
    34.01362, 30.8263, 30.65885, 30.5353, 30.64653, 30.82378, 31.51835,
    32.2942, 32.52289, 31.48866, 30.11888, 29.21234, 28.13532, 27.60697,
    27.38679, 27.1793, 27.09031, 27.21216, 27.72377, 27.81236, 27.28395,
    26.85345, 26.01127,
  17.51942, 17.54852, 17.57511, 17.59542, 17.58774, 17.57986, 17.5758,
    17.60159, 17.67225, 17.72164, 18.47816, 18.60351, 17.73919, 17.86926,
    17.98565, 17.69354, 17.61035, 17.65253, 17.67113, 18.12573, 18.3588,
    17.90627, 17.86628, 18.31015, 18.53326, 18.19283, 20.31577, 21.77198,
    19.17983, 18.08693,
  17.82634, 17.87228, 17.69601, 17.92702, 17.78548, 17.63183, 17.68118,
    17.74774, 17.83814, 17.97724, 18.33351, 18.82249, 19.05274, 18.4584,
    18.19825, 18.20988, 17.76249, 17.7886, 18.15165, 18.57899, 18.51504,
    18.02378, 18.02013, 18.71351, 22.06203, 22.48819, 21.12912, 24.07307,
    20.03704, 18.6303,
  17.77694, 17.79921, 17.7692, 17.82009, 17.7526, 17.69218, 17.71595,
    17.80642, 17.89963, 17.94927, 18.03423, 18.40327, 18.6635, 19.06139,
    19.14122, 18.35352, 18.26165, 18.55708, 18.51916, 18.69306, 19.39768,
    20.5607, 21.55154, 21.14091, 25.65632, 28.38108, 23.62822, 23.97989,
    20.09819, 19.23748,
  17.78355, 17.78997, 17.95297, 18.10168, 18.3418, 18.74856, 18.78809,
    18.56528, 18.60017, 18.87327, 18.92349, 19.17751, 19.01219, 18.67222,
    19.52098, 20.30776, 19.68155, 18.75583, 18.87713, 19.18788, 21.57217,
    23.0221, 22.08247, 26.60166, 28.54406, 25.46306, 26.49046, 23.50763,
    20.04488, 18.60344,
  18.27081, 17.99225, 18.23174, 18.55131, 18.87616, 19.06384, 19.03974,
    18.89447, 19.39691, 19.78752, 19.5362, 19.38337, 19.1935, 19.42789,
    20.11584, 20.50214, 19.6276, 18.99866, 19.4195, 23.89785, 25.7689,
    21.27702, 21.16101, 23.20917, 24.7493, 24.29275, 23.41659, 23.45582,
    24.08059, 20.18324,
  18.35553, 18.42332, 19.10027, 20.0518, 20.0006, 19.57245, 19.64515,
    19.41073, 19.09589, 19.16771, 19.153, 20.72999, 22.74832, 22.90392,
    22.30437, 28.6766, 35.62302, 28.11398, 22.56594, 24.63754, 23.22378,
    20.00601, 20.48556, 21.12341, 23.60198, 23.22093, 25.17447, 37.08864,
    33.92646, 19.65693,
  18.79766, 19.12264, 19.87827, 20.74858, 20.78946, 20.49033, 21.19679,
    22.64594, 22.95261, 22.80135, 23.38053, 23.25042, 22.4178, 22.45488,
    27.43981, 34.89509, 32.61755, 25.10949, 22.53887, 22.26058, 20.82453,
    19.90096, 20.44007, 22.71525, 24.22729, 21.46161, 30.15377, 45.5431,
    34.10075, 18.26354,
  19.6658, 20.04817, 20.97003, 21.96218, 21.86723, 23.74445, 26.07206,
    24.30823, 22.81447, 22.8442, 22.71198, 21.84597, 20.93657, 21.14396,
    23.45667, 25.36025, 23.98095, 22.46986, 21.04049, 20.78717, 20.20623,
    19.88481, 21.24253, 23.66006, 23.3267, 21.46133, 33.69839, 39.83272,
    24.37238, 18.45537,
  22.34332, 22.63166, 23.73768, 24.10225, 24.53869, 26.3988, 25.7145,
    24.04422, 23.74112, 23.487, 22.59087, 21.51724, 20.93756, 24.01565,
    25.99363, 22.77705, 22.70347, 24.28697, 24.10954, 21.93949, 20.05762,
    21.43585, 25.48686, 26.32026, 22.86094, 23.23839, 30.02121, 28.98371,
    20.38015, 18.50469,
  26.49905, 28.14788, 29.68148, 31.2164, 31.27241, 28.28645, 24.53725,
    24.20428, 23.43734, 22.42872, 22.989, 25.97246, 27.39991, 27.21517,
    25.80355, 25.73041, 26.43756, 26.89434, 25.3499, 23.66903, 23.68018,
    24.38938, 25.62629, 24.20482, 28.68407, 38.05247, 32.12033, 21.50758,
    18.98679, 17.79089,
  38.3725, 41.49509, 38.54604, 34.49842, 33.09316, 31.50524, 27.7685,
    29.2944, 30.34694, 36.9851, 40.73611, 27.84664, 24.37491, 23.9507,
    23.34591, 24.29105, 25.48742, 25.25915, 23.92339, 23.61225, 25.97317,
    25.79026, 23.05806, 21.14029, 25.1198, 29.49247, 24.05651, 18.55409,
    18.09967, 17.61495,
  53.9302, 43.28003, 44.95856, 46.15662, 44.56019, 38.84239, 41.70478,
    39.05254, 32.14162, 36.58821, 36.23832, 23.00502, 23.81411, 24.68653,
    23.03135, 23.56648, 23.05989, 22.78794, 22.2358, 22.71429, 25.58976,
    24.75397, 20.73205, 23.77685, 25.72842, 20.42605, 18.10214, 18.40438,
    18.28561, 17.77893,
  62.20144, 57.6645, 73.20556, 78.8665, 79.32314, 71.03493, 54.97026,
    36.67347, 33.94034, 32.08509, 28.84972, 21.48006, 25.70781, 28.23166,
    24.22113, 23.43417, 23.47875, 22.71043, 22.0139, 24.19188, 25.95875,
    23.04101, 20.36604, 25.2421, 26.75871, 19.62161, 18.21063, 18.54177,
    18.77187, 18.05549,
  69.03631, 93.45525, 95.46761, 92.5271, 82.25838, 70.50218, 59.15094,
    53.13976, 44.21487, 38.91703, 44.38285, 42.46486, 44.91661, 44.1098,
    37.95713, 29.85854, 23.93841, 25.27527, 26.62472, 27.81706, 25.31149,
    23.99179, 25.7341, 23.12594, 20.6733, 18.75373, 18.2584, 18.1466,
    18.48832, 18.02539,
  52.77599, 61.58028, 59.8698, 57.49862, 50.69483, 52.79554, 69.19102,
    66.87904, 57.2083, 56.86914, 55.17284, 42.5117, 33.14218, 38.02434,
    40.04926, 27.94857, 27.16968, 27.51725, 30.38538, 31.50792, 27.6315,
    24.90639, 22.44674, 19.83267, 18.44642, 18.81137, 18.34999, 18.01555,
    18.01468, 17.78795,
  41.60337, 41.42986, 40.70168, 38.81153, 37.40464, 41.66547, 48.65968,
    46.44428, 42.91016, 41.65869, 38.53981, 30.17487, 25.16626, 29.2516,
    29.38286, 26.73263, 28.54575, 27.14461, 28.20655, 28.12311, 23.31162,
    20.95062, 18.89696, 18.74259, 18.95062, 18.76657, 18.39884, 18.10236,
    17.95946, 17.71745,
  39.0098, 37.54723, 35.76631, 34.70635, 35.13194, 36.05196, 36.40991,
    35.96278, 34.45158, 32.11385, 27.43588, 26.22999, 29.30474, 27.94461,
    26.69427, 27.03955, 27.10787, 25.16128, 26.28926, 25.28761, 19.67143,
    19.54206, 19.24457, 18.92449, 18.78056, 18.76499, 18.34474, 17.92274,
    17.87925, 17.71453,
  35.14665, 34.06282, 32.94866, 33.23632, 33.53235, 34.11706, 34.26344,
    33.73983, 32.29337, 28.43129, 26.65651, 29.15647, 29.83963, 29.14179,
    30.56696, 28.85246, 25.06627, 22.7803, 25.22394, 24.15294, 19.61756,
    19.91404, 19.68407, 19.2095, 18.46486, 18.50504, 18.2371, 17.76521,
    17.73591, 17.64095,
  34.30439, 34.11474, 32.75824, 32.27412, 32.42056, 32.21096, 31.91544,
    31.08507, 28.93002, 26.52033, 28.00306, 28.58157, 25.18207, 25.79294,
    26.74688, 25.60882, 24.92821, 25.31267, 27.5701, 26.47955, 22.43711,
    20.83794, 19.95704, 19.38877, 18.39616, 18.21428, 18.09066, 17.76628,
    17.69269, 17.6209,
  34.56334, 34.50606, 32.9205, 31.4221, 31.29468, 30.91019, 30.31638,
    29.34409, 27.90161, 28.63817, 29.26575, 25.42637, 22.83347, 22.89028,
    22.71607, 22.03813, 23.18991, 25.1404, 26.85959, 27.37982, 25.53886,
    22.6089, 20.14554, 19.49982, 18.74564, 18.25153, 18.02278, 17.7813,
    17.68819, 17.62034,
  34.14234, 34.12164, 32.34879, 30.78657, 30.35665, 30.16172, 29.78837,
    29.08209, 28.70981, 29.8171, 27.49322, 22.54977, 22.19709, 22.26282,
    21.78908, 21.09163, 21.41841, 22.19743, 23.33941, 23.91091, 23.84933,
    23.30248, 21.68204, 20.11591, 19.13483, 18.50323, 18.03134, 17.78816,
    17.69743, 17.61814,
  34.59841, 33.49821, 31.77994, 30.68111, 30.34765, 29.92518, 29.87458,
    29.35877, 29.7421, 29.27332, 24.7255, 21.19931, 21.41459, 21.43932,
    21.16724, 20.98011, 20.72751, 20.64223, 20.92726, 20.83846, 21.88318,
    22.38482, 21.91408, 22.28541, 20.92846, 19.01856, 18.15107, 17.89268,
    17.72626, 17.63125,
  34.26542, 33.35435, 31.40967, 30.37723, 30.95011, 31.44412, 31.25268,
    30.01335, 29.88456, 27.63596, 22.66164, 20.7992, 20.82333, 20.87323,
    20.61847, 21.02558, 20.91162, 20.02532, 19.72972, 19.63124, 20.89835,
    21.08637, 20.17399, 21.89102, 22.26213, 19.92794, 18.39735, 18.27666,
    17.97757, 17.66721,
  33.67348, 32.92092, 32.0133, 31.81553, 32.22711, 32.36937, 32.5734,
    31.95586, 31.48963, 27.28301, 22.12026, 21.33684, 21.44134, 21.74939,
    21.62316, 21.64479, 21.66307, 20.80424, 19.82386, 19.75355, 20.13246,
    19.99884, 19.61333, 20.07763, 21.24617, 21.40596, 19.82032, 18.60769,
    18.32887, 17.80509,
  33.44197, 34.21732, 32.22881, 31.68292, 32.22329, 32.18518, 31.61088,
    31.2348, 31.64585, 27.54113, 22.24548, 21.67455, 21.84421, 22.09923,
    22.10486, 22.14816, 21.83639, 21.3984, 20.46743, 19.63657, 19.77474,
    19.89925, 19.8211, 19.35524, 19.25341, 20.53522, 20.52831, 19.24075,
    19.07859, 18.17852,
  33.88256, 35.9992, 34.65751, 33.09184, 32.0788, 31.12948, 31.63943, 32.286,
    30.77193, 26.46664, 22.78712, 22.18005, 22.44235, 22.14558, 21.63571,
    21.72268, 21.40545, 21.16749, 20.65906, 19.76009, 20.02107, 20.1875,
    19.45656, 18.90082, 18.82716, 19.438, 20.70174, 19.94516, 19.10007,
    18.15433,
  35.05345, 37.10142, 34.48838, 32.39738, 31.35273, 30.37185, 31.70633,
    32.3452, 29.10981, 25.05964, 23.13716, 22.50183, 22.24717, 21.78685,
    21.4617, 21.30212, 20.9525, 20.84583, 20.44476, 19.64872, 20.12794,
    21.2808, 21.39234, 20.54057, 20.23817, 20.41253, 22.13995, 21.83858,
    19.08894, 17.66768,
  34.83026, 35.38102, 32.99729, 31.94601, 32.16046, 31.69986, 32.48874,
    31.20365, 27.07329, 24.48421, 22.87435, 22.1488, 21.74088, 21.53347,
    21.8121, 21.5739, 20.87381, 20.60976, 20.79842, 21.00707, 21.936,
    22.31598, 21.72791, 20.8954, 20.77724, 20.90383, 21.36808, 23.2021,
    21.6257, 18.28991,
  32.31776, 31.41369, 31.6387, 32.82813, 33.84649, 34.92922, 33.909,
    29.87572, 26.34172, 24.39602, 22.07788, 20.69279, 20.37991, 20.71874,
    21.47585, 21.8489, 21.83625, 22.11355, 21.63462, 20.99224, 21.21827,
    20.92653, 20.01526, 19.49468, 19.74047, 20.18804, 20.31024, 20.54897,
    21.13394, 18.8926,
  30.78045, 30.92099, 31.27686, 31.56593, 32.07207, 34.53621, 34.76297,
    29.72262, 25.80135, 24.27442, 22.82774, 22.19124, 22.25526, 22.61122,
    22.97512, 23.14127, 22.27147, 21.23516, 20.6871, 19.87337, 19.40306,
    19.26875, 19.03169, 18.88507, 18.9886, 19.51444, 19.71368, 19.18616,
    18.7507, 17.91575,
  13.06113, 13.09061, 13.1148, 13.12583, 13.12719, 13.1169, 13.11665,
    13.13253, 13.17135, 13.2059, 13.92126, 13.97996, 13.21932, 13.40364,
    13.5077, 13.21796, 13.1549, 13.18093, 13.17654, 13.61712, 13.8098,
    13.401, 13.35307, 13.71649, 13.83317, 13.4729, 15.53684, 16.93214,
    14.76517, 13.64433,
  13.37471, 13.38717, 13.23204, 13.43463, 13.30025, 13.16654, 13.19532,
    13.2391, 13.30892, 13.44205, 13.8417, 14.32405, 14.47932, 13.92308,
    13.72314, 13.694, 13.28403, 13.3, 13.64235, 14.07672, 13.99296, 13.43094,
    13.36095, 13.91549, 16.90547, 17.20361, 16.60447, 19.38977, 15.70342,
    14.19066,
  13.32138, 13.33129, 13.29744, 13.34049, 13.26322, 13.19399, 13.20116,
    13.27382, 13.36276, 13.41725, 13.50378, 13.88887, 14.15224, 14.45984,
    14.48797, 13.77318, 13.68484, 13.92538, 13.87242, 13.97724, 14.48201,
    15.40636, 16.22579, 15.71506, 20.05404, 22.59642, 18.82312, 19.29716,
    15.6154, 14.71554,
  13.27632, 13.26013, 13.44441, 13.57408, 13.74956, 14.11399, 14.11733,
    13.87724, 13.92047, 14.1839, 14.24703, 14.5031, 14.28222, 14.02682,
    14.78528, 15.42956, 14.83466, 13.92945, 13.88361, 14.00625, 16.18949,
    17.53326, 16.78301, 20.83885, 22.56988, 20.52098, 21.57743, 18.78309,
    15.50326, 14.13794,
  13.64927, 13.40279, 13.62535, 13.91167, 14.22072, 14.3481, 14.25585,
    14.0925, 14.65771, 15.15637, 15.00131, 14.74176, 14.36164, 14.46494,
    15.11301, 15.41565, 14.3911, 13.72673, 14.05413, 18.25893, 19.90242,
    16.06623, 16.00357, 18.19345, 19.67775, 19.19374, 18.56815, 18.70752,
    18.99033, 15.32765,
  13.59862, 13.6024, 14.26324, 15.21737, 15.24697, 14.72892, 14.66305,
    14.47106, 14.25771, 14.37714, 14.2519, 15.53337, 17.14903, 17.32204,
    16.60633, 21.96647, 27.63766, 21.25639, 16.77123, 19.18482, 17.98847,
    14.92747, 15.48311, 16.10722, 18.41096, 18.01568, 19.86831, 30.28227,
    27.43791, 14.93175,
  13.66019, 13.93803, 14.70091, 15.65186, 15.79135, 15.29743, 15.70586,
    16.99628, 17.30962, 17.22668, 17.69484, 17.48361, 16.7783, 16.67254,
    20.98156, 27.77148, 26.21286, 19.36082, 17.12654, 17.04807, 15.7468,
    14.9189, 15.36843, 17.30625, 18.6997, 16.47031, 24.36808, 38.38639,
    28.57819, 13.68942,
  13.81689, 14.13163, 15.00001, 15.88721, 15.7646, 17.38696, 19.28257,
    17.78964, 16.74145, 16.93217, 16.97607, 16.09934, 15.18636, 15.31592,
    17.8254, 19.90948, 18.54071, 17.01707, 15.90949, 15.70376, 15.18647,
    14.91543, 16.00534, 18.07946, 17.91774, 15.98911, 28.24629, 34.53438,
    19.59468, 13.88736,
  15.1377, 15.28654, 16.3119, 16.51875, 16.91282, 18.89725, 18.41157,
    16.78881, 16.81054, 16.98901, 16.42618, 15.511, 15.10286, 18.1144,
    19.93604, 17.28809, 17.24245, 18.51711, 18.3342, 16.49276, 14.86684,
    15.90402, 19.4067, 20.26141, 17.37611, 17.30217, 24.07457, 23.76397,
    15.56268, 13.97134,
  17.2825, 18.51833, 20.00909, 21.22327, 21.57309, 19.2364, 16.21981,
    16.05097, 15.87455, 15.34524, 16.36846, 19.40848, 20.63806, 20.69945,
    19.99538, 19.89012, 20.44984, 20.84265, 19.78977, 18.56414, 18.47292,
    19.30628, 20.53892, 19.11655, 23.01082, 31.61766, 26.48851, 16.85087,
    14.51476, 13.31968,
  26.00055, 28.80362, 26.73445, 23.05326, 22.43591, 21.56846, 18.68198,
    20.36509, 21.8235, 28.05589, 31.43807, 21.40503, 18.64861, 18.32235,
    17.86168, 18.87136, 20.14141, 20.10403, 19.02249, 18.88944, 21.23723,
    21.28118, 18.67643, 16.58021, 20.52611, 25.26007, 20.09382, 14.22979,
    13.60558, 13.13735,
  39.23114, 29.93986, 31.38857, 32.40958, 31.37783, 27.34612, 30.44341,
    28.73306, 23.62558, 28.42056, 28.50973, 17.35939, 18.08585, 19.09788,
    17.89824, 18.43637, 18.11255, 18.02813, 17.65001, 18.16164, 21.05752,
    20.30207, 16.31159, 19.33557, 21.50875, 16.24749, 13.67758, 13.84466,
    13.7354, 13.28225,
  45.01112, 40.89025, 56.65026, 62.50876, 63.52487, 56.63286, 42.8889,
    27.39909, 25.52993, 24.69945, 21.96922, 15.70368, 20.13329, 22.58077,
    19.08353, 18.43874, 18.71436, 18.05712, 17.4275, 19.70768, 21.58711,
    18.62753, 15.92737, 21.05918, 22.88886, 15.28197, 13.68623, 13.98402,
    14.1777, 13.55417,
  53.28407, 76.71262, 79.1708, 76.6994, 68.00855, 58.31227, 48.46718,
    42.02578, 34.33221, 29.55529, 34.76289, 34.81489, 38.43147, 37.95697,
    31.79136, 24.48955, 19.17313, 20.43192, 21.66313, 22.87581, 20.75464,
    19.55052, 21.35771, 19.02183, 16.49062, 14.21714, 13.71692, 13.62026,
    13.95829, 13.54365,
  40.54403, 49.60041, 48.87003, 47.21598, 41.08727, 42.9206, 57.22338,
    54.79344, 44.53899, 44.41972, 45.51066, 35.54523, 27.80401, 32.7241,
    34.61247, 23.10378, 22.17237, 22.30533, 24.10295, 25.54796, 23.29657,
    20.78476, 18.52426, 15.64936, 13.81773, 14.18437, 13.78807, 13.49723,
    13.50804, 13.30833,
  30.07085, 30.43792, 30.54934, 29.5392, 28.19691, 32.53325, 39.86151,
    37.35563, 33.95752, 34.0914, 32.00224, 24.57781, 19.87567, 24.32956,
    24.80026, 21.77418, 23.53022, 21.96014, 22.09124, 22.50959, 19.23663,
    16.92464, 14.61497, 14.35992, 14.44009, 14.16994, 13.82942, 13.5843,
    13.44485, 13.23282,
  28.1892, 27.43818, 26.25067, 25.32694, 25.48046, 26.478, 27.17912,
    26.98969, 26.54483, 25.59197, 21.79282, 21.2573, 23.89716, 22.52469,
    21.78185, 21.95751, 22.13593, 20.0909, 20.51493, 19.90017, 15.19935,
    15.04239, 14.74877, 14.49891, 14.31572, 14.21452, 13.79314, 13.41752,
    13.38804, 13.23625,
  25.32845, 24.4947, 23.37337, 23.48973, 23.81881, 24.548, 25.11729,
    25.35751, 24.8752, 22.4191, 21.34099, 24.18334, 25.08889, 24.00376,
    25.22449, 23.69853, 20.34997, 18.0335, 19.8542, 18.90425, 14.89936,
    15.13762, 14.97843, 14.67392, 14.00243, 13.9883, 13.7476, 13.27996,
    13.25105, 13.17221,
  24.78076, 24.51261, 23.01819, 22.58195, 22.91484, 23.14376, 23.44427,
    23.36581, 22.22989, 20.90972, 22.87173, 23.98083, 20.97066, 21.31458,
    22.10829, 20.98195, 20.01901, 19.97468, 21.56248, 20.36487, 17.14359,
    15.94004, 15.16727, 14.79782, 13.90915, 13.71105, 13.60437, 13.29262,
    13.22388, 13.15057,
  24.9964, 24.95345, 23.4162, 22.09124, 22.23535, 22.1969, 22.10127,
    21.86562, 21.31694, 22.81474, 24.19393, 21.11439, 18.60502, 18.42654,
    18.15868, 17.58894, 18.41263, 19.95073, 20.98413, 21.13208, 20.03728,
    17.72656, 15.36834, 14.85595, 14.19439, 13.73468, 13.53429, 13.30185,
    13.22, 13.1528,
  24.57595, 24.70262, 23.19237, 21.89046, 21.69507, 21.67635, 21.63308,
    21.6041, 22.09724, 24.0911, 22.89948, 18.52443, 18.05407, 17.76759,
    16.99857, 16.34596, 16.59891, 17.29901, 18.0119, 18.43141, 18.89609,
    18.60079, 16.8165, 15.46377, 14.62763, 13.98457, 13.53732, 13.30387,
    13.22498, 13.15409,
  25.14449, 24.41663, 22.92134, 22.05728, 21.84135, 21.46559, 21.75265,
    21.97294, 23.15986, 23.889, 20.58713, 17.14032, 17.11564, 16.82009,
    16.29757, 16.06866, 15.89383, 15.83399, 16.18211, 16.22282, 17.33417,
    17.68703, 16.77717, 17.17224, 16.1007, 14.43803, 13.66349, 13.41245,
    13.24241, 13.15483,
  25.15582, 24.56937, 22.79101, 21.8763, 22.47697, 22.96722, 23.20012,
    22.68679, 23.32762, 22.5338, 18.63316, 16.57649, 16.32656, 16.1072,
    15.72627, 16.09994, 16.06601, 15.3461, 15.22098, 15.18149, 16.42447,
    16.4528, 15.16679, 16.7456, 17.24671, 15.27782, 13.89183, 13.78011,
    13.49199, 13.19053,
  24.79222, 24.40751, 23.44107, 23.27147, 23.92272, 24.21852, 24.74844,
    24.72193, 24.92844, 21.95607, 17.77619, 16.88717, 16.7052, 16.78526,
    16.51222, 16.58521, 16.70788, 15.98079, 15.20337, 15.2312, 15.57589,
    15.32831, 14.7784, 15.16063, 16.23251, 16.5647, 15.23388, 14.07951,
    13.8118, 13.31467,
  24.84083, 25.68478, 23.87222, 23.46592, 24.23725, 24.36802, 24.06982,
    24.02711, 24.98806, 22.04835, 17.68818, 17.09921, 16.94339, 17.08978,
    17.05492, 17.0535, 16.80766, 16.42098, 15.72362, 15.20567, 15.19614,
    15.14459, 15.06354, 14.66705, 14.63669, 15.94885, 15.99498, 14.70495,
    14.56238, 13.70664,
  25.36967, 27.57812, 26.29499, 24.76187, 24.19922, 23.49688, 23.86098,
    24.6172, 23.82569, 21.00671, 18.18236, 17.53419, 17.46621, 17.20351,
    16.71554, 16.74766, 16.44723, 16.21934, 15.97512, 15.38602, 15.40179,
    15.41786, 14.82398, 14.37597, 14.323, 14.91348, 16.10263, 15.36423,
    14.60203, 13.71136,
  26.66815, 29.02217, 26.6217, 24.44144, 23.50481, 22.45975, 23.81254,
    24.65627, 22.26464, 19.65779, 18.64009, 18.02402, 17.49405, 16.98892,
    16.59187, 16.41431, 16.10486, 16.04965, 15.90504, 15.32632, 15.46324,
    16.2876, 16.36647, 15.82805, 15.71408, 15.81998, 17.54113, 17.21802,
    14.56898, 13.23439,
  26.94173, 27.93613, 25.19964, 23.71686, 23.80682, 23.1902, 23.96081,
    23.37016, 20.57858, 19.25211, 18.54439, 17.79482, 17.00802, 16.70144,
    16.93906, 16.73764, 16.09156, 15.85028, 16.2365, 16.65825, 17.09177,
    17.16806, 16.77725, 16.31916, 16.36917, 16.35966, 16.84737, 18.60123,
    17.07665, 13.8297,
  24.73008, 23.71904, 23.58932, 24.74834, 25.33881, 25.57148, 24.86982,
    22.14554, 19.96381, 19.23117, 17.71721, 16.44057, 15.94577, 16.02415,
    16.6493, 16.98585, 16.89558, 17.14915, 16.98079, 16.65289, 16.72025,
    16.37956, 15.5387, 15.09231, 15.35572, 15.70173, 15.79313, 16.1397,
    16.72878, 14.44014,
  23.07144, 22.8901, 23.25663, 23.8009, 24.09357, 25.62794, 25.71925,
    22.13821, 19.51213, 18.99104, 18.05217, 17.55245, 17.72479, 17.75239,
    17.75456, 17.99003, 17.34425, 16.49592, 16.11575, 15.43064, 14.98072,
    14.90788, 14.64803, 14.47475, 14.56486, 15.06823, 15.28059, 14.72934,
    14.31425, 13.48037,
  9.742868, 9.753646, 9.779836, 9.799862, 9.795651, 9.788032, 9.79183,
    9.801814, 9.832011, 9.842418, 10.50015, 10.59224, 9.876934, 10.04697,
    10.16899, 9.903901, 9.825338, 9.840915, 9.828599, 10.21264, 10.41325,
    10.06285, 10.00779, 10.32585, 10.43369, 10.09063, 12.06617, 13.51467,
    11.5126, 10.39395,
  10.0093, 10.02084, 9.870502, 10.07735, 9.976194, 9.836881, 9.852607,
    9.890082, 9.941807, 10.06277, 10.50844, 10.95671, 11.09726, 10.61784,
    10.39866, 10.3696, 9.953344, 9.94681, 10.26421, 10.70305, 10.65753,
    10.09807, 9.981375, 10.47346, 13.45228, 13.87404, 13.48325, 16.55109,
    12.66485, 11.01058,
  10.00634, 10.00627, 9.949656, 10.01777, 9.938506, 9.839768, 9.838534,
    9.907216, 9.997929, 10.06669, 10.14345, 10.52997, 10.86519, 11.10774,
    11.08517, 10.41313, 10.2887, 10.52343, 10.48482, 10.56988, 10.97012,
    11.76064, 12.54762, 11.97331, 16.52557, 19.59373, 15.81823, 16.6264,
    12.5714, 11.59375,
  9.956321, 9.913913, 10.06711, 10.16451, 10.29067, 10.63138, 10.65408,
    10.42796, 10.46386, 10.73706, 10.84427, 11.08409, 10.85809, 10.64315,
    11.34142, 11.83416, 11.33468, 10.52759, 10.36797, 10.33646, 12.34536,
    13.77404, 13.09871, 17.08116, 19.14634, 17.41611, 18.78261, 16.00397,
    12.46476, 10.99901,
  10.28058, 10.00246, 10.18643, 10.42139, 10.7181, 10.91684, 10.82327,
    10.60172, 11.13761, 11.77264, 11.73636, 11.38828, 10.89156, 10.94989,
    11.63537, 11.89636, 10.77544, 10.04213, 10.2663, 14.07983, 15.89803,
    12.52258, 12.41559, 14.87711, 16.39966, 15.79589, 15.63262, 15.73701,
    15.76079, 12.01041,
  10.19059, 10.10321, 10.65128, 11.5445, 11.70792, 11.26545, 11.11904,
    10.94855, 10.8346, 10.99977, 10.85276, 11.87899, 13.33531, 13.55088,
    12.6828, 17.31085, 22.59785, 16.92484, 12.78419, 15.37439, 14.51028,
    11.46363, 12.07476, 12.64002, 14.86861, 14.66374, 16.07246, 26.70751,
    24.66603, 11.70586,
  10.14233, 10.37586, 11.09817, 12.06416, 12.34432, 11.80388, 11.95149,
    13.08319, 13.29354, 13.22819, 13.69541, 13.61918, 13.07534, 12.82133,
    16.7646, 23.79331, 22.71782, 15.73962, 13.55505, 13.60596, 12.34354,
    11.55205, 12.01902, 13.83284, 15.28541, 12.90669, 20.76576, 36.39014,
    26.75343, 10.35275,
  10.25592, 10.5574, 11.37687, 12.23226, 12.12613, 13.53019, 15.26451,
    13.90954, 12.91599, 13.13323, 13.29604, 12.44517, 11.39499, 11.36574,
    14.10407, 16.68829, 15.22012, 13.50963, 12.52913, 12.35172, 11.88067,
    11.60248, 12.58657, 14.65239, 14.6203, 12.33642, 25.10337, 33.11038,
    16.88572, 10.51959,
  11.37064, 11.47588, 12.42321, 12.59814, 12.90077, 15.09692, 14.80152,
    12.88302, 12.84531, 13.13437, 12.66236, 11.66226, 11.09664, 14.01115,
    15.99571, 13.59573, 13.72132, 15.15292, 14.89888, 13.10074, 11.51847,
    12.47836, 15.88099, 16.88768, 14.08633, 13.74699, 20.94089, 21.22136,
    12.04947, 10.67791,
  13.14541, 14.23576, 15.79472, 17.12291, 17.37968, 15.27623, 12.36001,
    12.03001, 11.87064, 11.34138, 12.17604, 15.0912, 16.56739, 16.94774,
    16.36553, 16.19073, 16.80013, 17.30198, 16.41465, 15.26826, 15.09495,
    15.99267, 17.4147, 16.06302, 19.61585, 28.36071, 23.64565, 13.72168,
    11.2416, 10.01281,
  20.28116, 23.13633, 21.55705, 18.25525, 17.73561, 17.17261, 14.36693,
    15.69584, 16.81093, 22.65169, 26.37823, 17.52517, 15.28034, 15.04175,
    14.52748, 15.55623, 16.90707, 16.90086, 15.75448, 15.58261, 17.92748,
    18.09398, 15.56979, 13.39049, 17.58132, 22.97358, 17.68636, 11.02483,
    10.28646, 9.794168,
  32.37573, 23.97198, 25.49256, 26.29407, 25.25485, 21.18663, 24.61353,
    23.51761, 18.50099, 23.52199, 24.51089, 13.98354, 14.72625, 15.82389,
    14.70415, 15.22598, 14.84947, 14.76596, 14.3731, 14.85561, 17.76378,
    17.1191, 13.0346, 15.99651, 18.61941, 13.39408, 10.46511, 10.51071,
    10.40569, 9.959326,
  40.38275, 33.94253, 45.90147, 52.11535, 54.4315, 50.21439, 37.97661,
    21.651, 20.53879, 20.35678, 18.06989, 12.23765, 16.83792, 19.46845,
    15.85482, 15.02609, 15.2477, 14.58991, 14.05227, 16.55726, 18.52823,
    15.36479, 12.59358, 18.09232, 20.45953, 12.17304, 10.38318, 10.66968,
    10.86857, 10.2629,
  47.79347, 68.87141, 72.01164, 74.02051, 70.41102, 59.31107, 41.71638,
    36.66531, 29.30298, 24.63005, 30.00368, 30.52833, 34.09411, 33.99798,
    28.04196, 21.10419, 15.63475, 16.99496, 18.39333, 19.82974, 17.72872,
    16.50331, 18.76884, 16.39584, 13.71735, 10.93167, 10.41979, 10.31253,
    10.67349, 10.28117,
  34.18325, 43.0745, 43.96117, 45.41515, 40.87145, 39.94016, 50.93957,
    50.46077, 39.95686, 40.06261, 41.80414, 32.21741, 24.53203, 29.2158,
    31.59693, 19.77773, 18.64146, 18.73578, 20.28018, 22.11553, 20.51639,
    18.20021, 16.11413, 12.77966, 10.44239, 10.84865, 10.48924, 10.20593,
    10.21448, 10.01148,
  23.66373, 24.2635, 25.17356, 24.78907, 22.91026, 27.01675, 35.03511,
    32.30933, 29.59434, 30.91504, 29.26007, 21.81537, 16.79876, 21.17716,
    21.71145, 18.42573, 20.303, 18.44335, 18.22752, 19.1586, 16.51682,
    14.22842, 11.60489, 11.19675, 11.15622, 10.84376, 10.5202, 10.29091,
    10.13764, 9.924438,
  22.24038, 21.90497, 21.13338, 20.17936, 20.09692, 21.24961, 22.05953,
    21.75283, 22.17637, 22.19104, 18.80536, 18.26037, 20.54441, 19.02832,
    18.48143, 18.86487, 19.15208, 16.84103, 16.99167, 16.80221, 12.18173,
    11.91114, 11.53809, 11.33127, 11.11135, 10.93188, 10.46931, 10.10145,
    10.05194, 9.915944,
  19.93192, 19.36926, 18.3185, 18.4035, 18.87818, 19.6567, 20.29868,
    20.92657, 20.83433, 18.9397, 17.88156, 20.72716, 21.97109, 20.77043,
    22.49807, 21.17085, 17.59743, 14.75294, 16.48661, 15.89004, 11.69025,
    11.76391, 11.55874, 11.40628, 10.78135, 10.70675, 10.46094, 9.946411,
    9.917671, 9.84607,
  19.68232, 19.46956, 18.00011, 17.60753, 18.04948, 18.46456, 18.92589,
    19.07456, 18.21354, 17.16981, 19.15504, 20.66166, 18.13188, 18.53343,
    19.61977, 18.47587, 17.21574, 16.47264, 17.97205, 17.02073, 13.57115,
    12.38107, 11.67539, 11.44364, 10.63536, 10.42097, 10.32226, 9.965331,
    9.89627, 9.826448,
  20.05046, 19.95089, 18.4779, 17.30398, 17.53032, 17.60521, 17.61597,
    17.42434, 16.9703, 18.6572, 20.60289, 18.25124, 15.97397, 15.77044,
    15.45289, 14.85785, 15.52014, 16.634, 17.33417, 17.56399, 16.38188,
    14.1284, 11.83416, 11.49863, 10.92837, 10.43451, 10.24563, 9.998249,
    9.89479, 9.831591,
  19.68051, 19.82513, 18.39936, 17.23449, 17.16306, 17.14459, 16.9696,
    16.84906, 17.45241, 19.95259, 19.75615, 16.06395, 15.69309, 15.1595,
    14.15172, 13.39319, 13.47367, 13.92492, 14.47786, 14.98769, 15.55601,
    15.14821, 13.16138, 12.14218, 11.41789, 10.74011, 10.26429, 9.994816,
    9.895041, 9.830645,
  20.2937, 19.64214, 18.25265, 17.49735, 17.30431, 16.75101, 16.80613,
    17.03822, 18.58885, 20.26032, 18.05578, 14.86702, 14.72758, 14.13035,
    13.32302, 12.89651, 12.60999, 12.48113, 12.88164, 12.96156, 14.09945,
    14.51703, 13.35192, 13.84886, 12.81125, 11.16597, 10.37719, 10.09514,
    9.90696, 9.83342,
  20.42152, 19.855, 18.1794, 17.25635, 17.65026, 17.8841, 18.1453, 17.94954,
    19.12818, 19.36311, 16.3482, 14.33402, 13.81159, 13.24361, 12.58272,
    12.78144, 12.80258, 12.14341, 12.00447, 11.94156, 13.25816, 13.40205,
    11.88133, 13.46836, 13.88989, 11.94581, 10.59482, 10.4998, 10.17356,
    9.858239,
  20.09463, 19.74112, 18.65487, 18.28537, 18.81552, 19.11694, 19.98904,
    20.47186, 21.09185, 18.78311, 15.3913, 14.53467, 14.01247, 13.73714,
    13.21273, 13.23346, 13.45318, 12.74994, 11.9229, 11.95798, 12.43075,
    12.17637, 11.51141, 11.90776, 12.87094, 13.14838, 11.90579, 10.81097,
    10.49702, 9.992791,
  19.97697, 20.44537, 18.81668, 18.44497, 19.36654, 19.92185, 20.0428,
    20.15544, 21.13376, 18.80717, 15.12014, 14.62547, 14.20981, 14.0282,
    13.79116, 13.78471, 13.5661, 13.15877, 12.44213, 11.99871, 11.99343,
    11.88817, 11.85398, 11.45543, 11.36181, 12.66954, 12.83114, 11.52165,
    11.27394, 10.43476,
  20.20148, 21.88974, 21.00288, 19.93502, 19.85753, 19.66753, 20.11378,
    20.74109, 19.94908, 17.77292, 15.39034, 14.92461, 14.68651, 14.15025,
    13.51365, 13.47607, 13.14157, 12.89948, 12.6729, 12.13471, 12.14879,
    12.16043, 11.58491, 11.09309, 11.01633, 11.66157, 12.94081, 12.21523,
    11.36798, 10.49993,
  21.36332, 23.29695, 21.73983, 20.24584, 19.60922, 18.74818, 20.18431,
    20.96262, 18.49665, 16.33239, 15.79012, 15.47253, 14.86074, 13.98149,
    13.29735, 12.9992, 12.72668, 12.67817, 12.55216, 12.02822, 12.12221,
    12.94127, 12.9858, 12.41954, 12.38971, 12.57005, 14.40641, 14.13025,
    11.37984, 9.999274,
  22.0974, 23.13588, 20.80656, 19.67639, 19.82741, 19.24878, 19.96252,
    19.43062, 16.70874, 15.8976, 15.82636, 15.38648, 14.40013, 13.59119,
    13.47376, 13.19207, 12.61983, 12.41368, 12.80244, 13.29267, 13.6116,
    13.70896, 13.39318, 12.94699, 13.08483, 13.17521, 13.78694, 15.48443,
    13.89031, 10.56369,
  20.67827, 19.9025, 19.73322, 20.95686, 21.34857, 21.13505, 20.47407,
    17.96733, 16.07793, 16.07042, 15.21732, 14.08025, 13.18289, 12.76974,
    13.11545, 13.41116, 13.36065, 13.65149, 13.5793, 13.36001, 13.42349,
    13.06544, 12.22927, 11.75702, 12.05954, 12.46731, 12.58549, 12.99843,
    13.57539, 11.2467,
  19.42876, 19.2424, 19.57895, 20.10776, 20.13109, 21.24868, 21.21622,
    17.898, 15.78591, 15.87745, 15.35136, 14.83139, 14.53776, 14.16909,
    14.15542, 14.49718, 13.94801, 13.14317, 12.7657, 12.13344, 11.68499,
    11.6312, 11.36908, 11.15968, 11.26591, 11.77375, 12.04706, 11.50699,
    11.07784, 10.22963,
  11.46094, 11.47458, 11.50139, 11.51808, 11.50708, 11.50891, 11.51537,
    11.52833, 11.55801, 11.55701, 12.21914, 12.40399, 11.60732, 11.73855,
    11.9097, 11.65888, 11.55953, 11.57161, 11.54923, 11.93598, 12.22148,
    11.85353, 11.76511, 12.08702, 12.17604, 11.78126, 13.7028, 15.40661,
    13.30693, 12.21249,
  11.71693, 11.77585, 11.5981, 11.81858, 11.70843, 11.56095, 11.58422,
    11.61089, 11.67176, 11.80636, 12.29089, 12.77794, 12.87564, 12.4077,
    12.17495, 12.20154, 11.71294, 11.6746, 12.00744, 12.52556, 12.52696,
    11.88925, 11.68991, 12.17218, 15.22701, 16.13799, 15.31769, 19.05075,
    14.64752, 12.92992,
  11.74245, 11.75787, 11.68108, 11.76876, 11.677, 11.55868, 11.55114,
    11.62426, 11.73512, 11.82219, 11.89668, 12.29088, 12.67454, 12.93746,
    12.96124, 12.23745, 12.04596, 12.33194, 12.30101, 12.39591, 12.76562,
    13.56202, 14.36947, 13.71958, 18.41939, 22.6461, 17.86606, 19.14176,
    14.54648, 13.60424,
  11.70252, 11.64358, 11.79143, 11.89698, 12.00782, 12.35686, 12.41083,
    12.17542, 12.17898, 12.4428, 12.58473, 12.85288, 12.67146, 12.42314,
    13.23401, 13.81058, 13.34251, 12.41347, 12.13929, 11.99341, 13.93847,
    15.65403, 14.81752, 18.92283, 21.8015, 19.71702, 21.36164, 18.41642,
    14.50443, 12.94715,
  12.09951, 11.72613, 11.91064, 12.13892, 12.45917, 12.72188, 12.64336,
    12.35455, 12.84125, 13.60554, 13.66621, 13.28201, 12.72557, 12.81111,
    13.61717, 13.94538, 12.71453, 11.73434, 11.83793, 15.64471, 18.06438,
    14.32397, 14.07112, 16.76988, 18.70749, 17.9814, 17.9709, 17.98301,
    18.00024, 14.02354,
  11.97892, 11.80953, 12.37194, 13.31066, 13.56143, 13.15093, 12.93871,
    12.72978, 12.61728, 12.84873, 12.70992, 13.68531, 15.31348, 15.62682,
    14.65353, 19.03395, 25.08209, 19.17962, 14.39419, 17.21445, 16.68573,
    13.17904, 13.81293, 14.53927, 16.92307, 17.00318, 17.76893, 29.4356,
    28.33546, 13.71467,
  11.83592, 12.05664, 12.83474, 13.90269, 14.27027, 13.69938, 13.70351,
    14.95746, 15.22528, 15.15213, 15.62602, 15.60347, 15.06175, 14.69362,
    18.96582, 27.20892, 26.06754, 17.86351, 15.32697, 15.51567, 14.21333,
    13.31149, 13.80741, 15.82166, 17.57467, 14.99199, 22.50077, 40.47664,
    31.46171, 12.22396,
  11.92242, 12.2458, 13.09105, 14.04808, 13.9318, 15.14741, 17.08554,
    15.9089, 14.80643, 15.09153, 15.32078, 14.44153, 13.16374, 13.01531,
    16.10185, 19.47233, 17.58344, 15.41262, 14.30774, 14.20063, 13.73793,
    13.40187, 14.44303, 16.69984, 16.81015, 14.09871, 27.95387, 38.78151,
    19.69803, 12.36462,
  13.0381, 13.14013, 14.10936, 14.33173, 14.49075, 16.91454, 16.85293,
    14.71596, 14.67276, 15.05325, 14.58391, 13.46603, 12.71218, 15.69479,
    18.18026, 15.60411, 15.5696, 17.23257, 17.0534, 15.1977, 13.30793,
    14.20589, 17.75175, 19.08852, 15.94497, 15.44134, 23.65263, 25.15936,
    13.91118, 12.55532,
  14.7856, 15.87183, 17.52516, 19.12536, 19.43657, 17.44271, 14.20201,
    13.82431, 13.7046, 13.14913, 13.70432, 16.83862, 18.54451, 19.04862,
    18.50699, 18.30113, 18.97647, 19.58227, 18.77132, 17.46803, 17.12835,
    18.01118, 19.60016, 18.04085, 21.80326, 32.15719, 27.34913, 16.06497,
    13.25971, 11.7936,
  21.84886, 25.20613, 23.96891, 20.56237, 19.85198, 19.50062, 16.3248,
    17.55161, 18.63116, 23.8275, 28.5615, 19.78373, 17.25502, 17.0432,
    16.48717, 17.66883, 19.32633, 19.32876, 18.0766, 17.63116, 20.14543,
    20.45173, 17.75902, 15.12029, 19.67617, 26.23829, 20.83208, 13.04698,
    12.13094, 11.52165,
  34.71744, 26.547, 27.5268, 27.98889, 27.24881, 22.08088, 25.8837, 25.67675,
    19.91185, 24.73647, 26.52311, 15.63443, 16.41432, 17.93287, 16.77335,
    17.5032, 17.13602, 17.03836, 16.50596, 16.90597, 19.98163, 19.46872,
    14.95975, 17.72415, 21.0133, 15.69765, 12.38988, 12.35663, 12.23369,
    11.72158,
  50.42933, 39.46067, 42.72319, 50.98824, 55.83082, 51.90241, 39.95139,
    22.17425, 21.44351, 21.40021, 19.48134, 13.30738, 18.32475, 21.60697,
    18.06563, 17.25415, 17.53172, 16.76546, 16.11711, 18.77444, 21.06107,
    17.55832, 14.45964, 20.04182, 23.47219, 14.40544, 12.21096, 12.50981,
    12.76915, 12.11237,
  51.65172, 68.13096, 66.03745, 72.47418, 71.25017, 60.83646, 42.38969,
    36.36778, 29.78803, 24.72292, 30.83833, 31.87905, 35.63443, 36.33807,
    30.68473, 24.37477, 17.88238, 19.38872, 20.83621, 22.44751, 20.24226,
    18.57506, 21.53935, 19.1502, 16.12429, 12.88953, 12.25074, 12.14507,
    12.5489, 12.13967,
  32.08086, 38.91895, 39.73252, 43.44214, 40.58069, 39.51172, 50.35695,
    50.04777, 39.56848, 40.03066, 43.62548, 33.4367, 26.01101, 31.47402,
    34.94624, 22.5309, 21.28233, 21.30529, 22.77221, 24.84739, 23.31754,
    20.79993, 18.81542, 15.29338, 12.33684, 12.7289, 12.34629, 12.02962,
    12.04389, 11.82735,
  20.73892, 21.14896, 22.91676, 23.04729, 21.25868, 24.84655, 32.99584,
    30.1162, 27.46436, 29.88156, 29.75284, 22.40497, 17.78125, 23.11146,
    24.33664, 20.84699, 23.09176, 21.1125, 20.57088, 21.7707, 19.05416,
    16.71032, 13.80295, 13.20143, 13.06814, 12.72124, 12.36072, 12.14523,
    11.97073, 11.7073,
  19.36367, 19.00761, 18.49933, 17.48638, 17.0935, 18.25629, 19.43488,
    19.0901, 19.48053, 20.45727, 17.85113, 18.02328, 21.55286, 20.6953,
    20.84167, 21.51677, 21.91437, 19.48732, 19.47911, 19.7262, 14.43601,
    14.09294, 13.57881, 13.34755, 13.05351, 12.77684, 12.29001, 11.90937,
    11.84365, 11.68358,
  16.95768, 16.3728, 15.23318, 15.15259, 15.55702, 16.55741, 17.44101,
    18.05819, 18.0252, 16.56145, 16.17073, 20.30752, 22.93135, 22.46164,
    25.41144, 24.23039, 20.26843, 17.13962, 19.02054, 18.78675, 13.86197,
    13.81893, 13.54684, 13.46877, 12.72988, 12.52379, 12.28171, 11.70246,
    11.66736, 11.58976,
  16.7634, 16.39139, 14.73533, 14.19009, 14.69925, 15.2634, 15.80485,
    15.95935, 15.2045, 14.35238, 17.19699, 20.20384, 18.62248, 20.17445,
    22.48927, 21.3996, 19.81582, 18.76183, 20.43351, 19.7448, 15.82348,
    14.42159, 13.66109, 13.46515, 12.53931, 12.23834, 12.1412, 11.72289,
    11.63054, 11.55209,
  17.06514, 16.69533, 15.16855, 13.88167, 14.18138, 14.30858, 14.34588,
    14.17231, 13.74355, 15.75152, 18.79824, 17.60354, 16.33195, 17.38086,
    17.89694, 17.40675, 18.04806, 19.09929, 19.63867, 19.96627, 18.71976,
    16.47554, 13.88434, 13.48993, 12.85319, 12.25449, 12.04291, 11.76815,
    11.6316, 11.56042,
  16.52174, 16.43208, 15.06609, 13.85013, 13.784, 13.82527, 13.65801,
    13.50584, 14.21086, 17.24542, 18.08067, 15.2556, 16.16856, 16.82837,
    16.38335, 15.70918, 15.78603, 16.18594, 16.61243, 17.25764, 18.07724,
    17.80099, 15.38141, 14.1707, 13.32531, 12.57819, 12.06435, 11.76096,
    11.63434, 11.5641,
  17.24721, 16.21747, 14.91463, 14.15498, 13.99201, 13.392, 13.46919,
    13.70511, 15.53151, 17.85509, 16.36771, 14.07221, 15.29925, 15.74095,
    15.40416, 15.0977, 14.7375, 14.53507, 15.0057, 15.20416, 16.57126,
    17.19083, 15.45806, 16.02917, 14.87214, 13.0819, 12.16992, 11.87401,
    11.65134, 11.56475,
  17.36331, 16.47783, 14.86147, 13.93507, 14.41979, 14.61823, 14.90996,
    14.80911, 16.30549, 17.05541, 14.5543, 13.57492, 14.31558, 14.69612,
    14.52126, 14.9092, 14.98643, 14.2701, 14.13623, 14.03128, 15.50134,
    15.86322, 13.76602, 15.57571, 16.11071, 13.97364, 12.38554, 12.28094,
    11.92402, 11.59369,
  17.08775, 16.48132, 15.44438, 15.06313, 15.67293, 16.03551, 17.1524,
    17.87829, 18.65163, 16.4957, 13.51355, 13.71842, 14.37819, 15.09135,
    15.17146, 15.43075, 15.74461, 14.98123, 13.99478, 13.98959, 14.51767,
    14.21689, 13.33051, 13.83271, 14.93409, 15.15439, 13.76541, 12.63411,
    12.28492, 11.74331,
  16.82774, 16.85308, 15.51573, 15.29962, 16.4344, 17.31916, 17.66558,
    17.78274, 18.75581, 16.57879, 13.17467, 13.72466, 14.53758, 15.39597,
    15.79487, 16.00973, 15.77656, 15.35023, 14.51386, 13.99745, 13.94113,
    13.76248, 13.7557, 13.3578, 13.23908, 14.62571, 14.8673, 13.47806,
    13.12657, 12.2662,
  16.94433, 17.8889, 17.5989, 17.0729, 17.22089, 17.38342, 17.98302,
    18.60848, 17.54141, 15.44833, 13.4091, 13.99282, 15.07436, 15.55836,
    15.41108, 15.53852, 15.23937, 15.00541, 14.7604, 14.15593, 14.06888,
    14.05811, 13.5212, 12.98116, 12.85133, 13.57237, 15.005, 14.30195,
    13.23026, 12.34448,
  18.07225, 19.22017, 18.46069, 17.59369, 17.11409, 16.45054, 18.1679,
    18.975, 16.08415, 13.79725, 13.79273, 14.59763, 15.35029, 15.43157,
    15.1625, 14.99581, 14.7558, 14.72609, 14.62425, 14.00663, 14.02514,
    14.88974, 15.02116, 14.37687, 14.3479, 14.57558, 16.49619, 16.29168,
    13.24878, 11.76855,
  19.20993, 19.85564, 17.6869, 17.17704, 17.4502, 16.92947, 17.84595,
    17.31801, 14.07145, 13.24471, 13.82762, 14.58545, 14.95199, 15.06599,
    15.40985, 15.26646, 14.63624, 14.39693, 14.78185, 15.25189, 15.60279,
    15.74874, 15.44407, 14.9731, 15.07496, 15.23138, 15.85231, 17.56726,
    16.0099, 12.42678,
  18.15978, 17.16948, 17.0168, 18.62665, 19.17719, 18.95647, 18.20658,
    15.45407, 13.17867, 13.38334, 13.18033, 13.19689, 13.58153, 14.13022,
    15.0027, 15.4409, 15.35823, 15.64288, 15.59877, 15.37781, 15.46363,
    15.03738, 14.16753, 13.67977, 13.97918, 14.44962, 14.56232, 14.95056,
    15.59787, 13.22087,
  17.45882, 17.20683, 17.6137, 18.17562, 18.39181, 19.3791, 19.0032,
    15.38232, 13.06623, 13.47438, 13.62918, 14.15411, 14.95832, 15.60842,
    16.10774, 16.52415, 15.98376, 15.1081, 14.68276, 14.06898, 13.59519,
    13.47381, 13.21435, 13.01524, 13.1383, 13.68322, 13.97354, 13.42462,
    12.94996, 12.03418,
  14.14452, 14.16541, 14.19128, 14.2087, 14.20079, 14.19608, 14.18643,
    14.20092, 14.22266, 14.21775, 14.85102, 15.12765, 14.29921, 14.44849,
    14.6767, 14.38824, 14.28079, 14.28885, 14.25489, 14.64675, 15.00906,
    14.62254, 14.49363, 14.83011, 14.91437, 14.4744, 16.38059, 18.53208,
    16.22727, 15.04656,
  14.37777, 14.47575, 14.27102, 14.51869, 14.40833, 14.22447, 14.23472,
    14.25515, 14.29681, 14.43155, 14.91671, 15.4422, 15.55841, 15.15334,
    14.91068, 14.9922, 14.44237, 14.37796, 14.72204, 15.29237, 15.35163,
    14.67368, 14.36002, 14.85186, 17.93669, 19.54139, 18.17256, 22.83666,
    17.77267, 15.88595,
  14.42778, 14.46062, 14.36928, 14.4825, 14.3749, 14.22654, 14.20539,
    14.27366, 14.37429, 14.47698, 14.56954, 14.96657, 15.41128, 15.73259,
    15.83145, 15.02878, 14.76339, 15.12381, 15.08677, 15.171, 15.54203,
    16.35904, 17.08526, 16.39126, 21.04188, 26.76662, 21.16054, 23.0355,
    17.64141, 16.63422,
  14.39843, 14.35022, 14.49888, 14.61835, 14.74051, 15.10446, 15.12493,
    14.85714, 14.84718, 15.10577, 15.29826, 15.64224, 15.51678, 15.18843,
    16.05225, 16.72297, 16.33582, 15.2444, 14.90715, 14.65288, 16.60489,
    18.6596, 17.51807, 21.79121, 25.77699, 23.08001, 25.40977, 22.16745,
    17.50739, 15.86372,
  14.87502, 14.44488, 14.65798, 14.86742, 15.20818, 15.49201, 15.37406,
    15.07025, 15.55308, 16.45372, 16.60739, 16.15722, 15.49135, 15.58509,
    16.46341, 16.84756, 15.55543, 14.39667, 14.47776, 18.35042, 21.60885,
    17.16771, 16.70009, 19.61664, 22.13855, 21.38995, 21.56228, 21.43106,
    21.37552, 17.02949,
  14.73417, 14.51495, 15.13225, 16.15085, 16.42077, 15.95842, 15.67326,
    15.44833, 15.35144, 15.66695, 15.51871, 16.47539, 18.40794, 18.70749,
    17.69082, 22.20366, 29.63939, 23.17643, 17.22472, 20.25119, 20.0268,
    15.82916, 16.45812, 17.35913, 19.9206, 20.55172, 20.32104, 32.39244,
    32.92353, 16.86561,
  14.55204, 14.7663, 15.62128, 16.84893, 17.314, 16.70601, 16.50428, 17.9228,
    18.32114, 18.22138, 18.69759, 18.84043, 18.27918, 17.74769, 22.05828,
    31.45892, 30.76143, 21.34603, 18.31126, 18.56129, 17.0821, 15.98715,
    16.56253, 18.79456, 20.89239, 18.25196, 24.4305, 44.61754, 38.29662,
    15.24011,
  14.62922, 14.98945, 15.92767, 17.02037, 16.9104, 18.14809, 20.42041,
    19.2193, 17.88408, 18.23516, 18.48887, 17.6476, 16.06872, 15.80718,
    19.06679, 23.1205, 20.84249, 18.36534, 17.18246, 17.00866, 16.54982,
    16.16174, 17.28268, 19.92982, 20.24456, 17.05228, 31.00037, 45.77264,
    24.46672, 15.36136,
  15.82881, 15.94342, 16.90473, 17.17791, 17.26672, 20.15986, 20.42839,
    17.77394, 17.66377, 18.17515, 17.72016, 16.38795, 15.41486, 18.39741,
    21.46053, 18.73266, 18.41189, 20.21935, 20.13935, 18.28323, 16.10469,
    17.05786, 20.86472, 22.77125, 19.18295, 18.456, 27.49335, 30.82726,
    17.11807, 15.5439,
  17.89433, 18.6584, 20.37545, 22.53035, 22.8968, 20.98503, 17.20345,
    16.70611, 16.56636, 16.01541, 16.42191, 19.86844, 21.67769, 22.23613,
    21.64763, 21.34994, 22.03734, 22.75619, 22.20042, 20.71681, 20.29026,
    21.16625, 22.97266, 21.53386, 24.93553, 36.81631, 33.02497, 19.81738,
    16.31988, 14.60375,
  23.53065, 27.53068, 27.33427, 23.53591, 22.89225, 22.85288, 19.32127,
    20.48082, 21.98856, 26.551, 32.47552, 23.64769, 20.45325, 20.11794,
    19.45159, 20.70064, 22.52779, 22.61891, 21.49147, 20.815, 23.63014,
    24.10581, 21.15862, 18.12751, 22.89587, 30.7035, 25.46925, 16.15678,
    15.00739, 14.23364,
  40.34215, 31.56175, 29.06646, 28.94849, 28.42169, 23.54238, 28.40514,
    29.29952, 23.14454, 28.08384, 30.74795, 18.61545, 19.18367, 20.90237,
    19.70031, 20.68846, 20.29746, 20.2103, 19.71714, 20.16145, 23.66162,
    23.29989, 18.08201, 20.77673, 25.29001, 19.71935, 15.52549, 15.18384,
    15.06391, 14.47581,
  54.57259, 38.54354, 42.74345, 50.58511, 55.67085, 52.59464, 43.37233,
    25.86276, 25.13193, 25.15339, 22.65426, 15.52754, 20.77457, 24.46236,
    21.2247, 20.39051, 20.79796, 19.99504, 19.14977, 22.11891, 25.01813,
    21.00257, 17.38948, 23.70962, 29.02803, 17.84266, 15.04106, 15.30727,
    15.58797, 14.92589,
  55.65081, 66.23906, 66.28335, 73.24683, 73.39591, 65.6515, 47.74613,
    40.4088, 34.02889, 28.5033, 33.97692, 34.50318, 39.71572, 41.37177,
    35.25035, 28.25458, 21.21322, 22.91908, 24.55783, 26.5084, 24.25141,
    21.78686, 25.83657, 23.73563, 20.34915, 15.89306, 15.05066, 14.93026,
    15.35072, 14.98343,
  35.2015, 40.58683, 42.9206, 49.23745, 48.41107, 45.88557, 55.33093,
    55.39233, 43.48417, 43.85419, 47.82841, 37.096, 29.73919, 36.16584,
    40.12047, 26.3996, 25.16591, 25.34482, 26.81796, 29.07055, 27.26844,
    24.74301, 23.2102, 19.29102, 15.22463, 15.57196, 15.15518, 14.83088,
    14.82882, 14.61164,
  23.09346, 24.24202, 27.65333, 29.26912, 27.2455, 29.18587, 37.26447,
    33.68298, 30.36998, 33.39552, 33.53243, 25.44215, 20.08648, 26.07229,
    27.98843, 24.29914, 27.22425, 25.23563, 24.23434, 25.72734, 22.80418,
    20.4985, 17.35, 16.35894, 15.95293, 15.55404, 15.14348, 14.92745,
    14.72588, 14.4499,
  21.65441, 22.10995, 22.23752, 20.98066, 19.85297, 20.90234, 22.33087,
    21.47429, 21.75431, 23.14729, 20.31159, 20.04534, 23.74579, 22.83445,
    23.56579, 24.87815, 25.97346, 23.43461, 23.15173, 24.12544, 18.02322,
    17.532, 16.67939, 16.30583, 15.96773, 15.63996, 15.09042, 14.69587,
    14.57661, 14.40259,
  19.21758, 19.01859, 17.68405, 17.2145, 17.42164, 18.53929, 19.44827,
    19.96969, 20.12834, 18.64975, 17.89242, 22.14683, 25.18443, 24.60239,
    28.82445, 28.15699, 24.16116, 20.66155, 22.81927, 23.32019, 17.29994,
    17.13256, 16.50384, 16.3955, 15.60895, 15.35517, 15.1286, 14.45951,
    14.39796, 14.30867,
  19.04716, 18.63545, 16.62948, 15.9062, 16.37585, 16.94034, 17.59068,
    17.85704, 17.23251, 16.15837, 18.7963, 22.08296, 20.45717, 22.30616,
    25.87128, 25.16352, 23.69015, 22.51861, 24.6307, 24.18566, 19.42188,
    17.73007, 16.59147, 16.37769, 15.36439, 15.01364, 14.92748, 14.46245,
    14.35964, 14.27592,
  19.32424, 18.68965, 16.92678, 15.47696, 15.75858, 15.93531, 16.11329,
    16.0659, 15.57385, 17.54109, 20.86466, 19.4491, 17.94151, 19.38759,
    20.60652, 20.58921, 21.69827, 23.25064, 23.88492, 24.13083, 22.44895,
    20.02658, 16.8921, 16.39173, 15.67033, 15.0212, 14.81187, 14.52556,
    14.35598, 14.28285,
  18.58832, 18.27024, 16.77019, 15.4401, 15.40147, 15.56856, 15.47172,
    15.25678, 15.94353, 19.25824, 20.42583, 17.03032, 17.84833, 18.77657,
    18.83215, 18.66632, 19.25109, 19.99145, 20.31688, 20.91959, 21.78315,
    21.61084, 18.5021, 17.11753, 16.1909, 15.4042, 14.84143, 14.51399,
    14.35492, 14.28811,
  19.35437, 17.97523, 16.64238, 15.83162, 15.76883, 15.16366, 15.19886,
    15.36391, 17.32759, 20.08617, 18.65032, 15.89248, 17.1605, 17.77811,
    17.86167, 18.05267, 18.08496, 17.86466, 18.28315, 18.48796, 19.92938,
    20.93048, 18.48355, 19.09217, 17.95971, 16.02357, 14.9403, 14.64649,
    14.36956, 14.27797,
  19.49358, 18.32089, 16.68067, 15.66289, 16.24782, 16.43758, 16.64371,
    16.49287, 18.22139, 19.41046, 16.72342, 15.524, 16.27082, 16.78492,
    16.92611, 17.74173, 18.1374, 17.43986, 17.24313, 17.09394, 18.69753,
    19.43515, 16.65567, 18.60548, 19.24208, 16.99942, 15.15106, 15.07186,
    14.67641, 14.31445,
  19.21856, 18.42746, 17.40479, 16.95392, 17.58815, 17.85413, 19.091,
    20.05527, 21.14377, 19.03801, 15.67353, 15.81957, 16.43491, 17.21157,
    17.52222, 18.19255, 18.85818, 18.19375, 17.0542, 17.02102, 17.76989,
    17.48987, 16.21586, 16.80904, 17.90567, 18.08652, 16.62782, 15.42046,
    15.04991, 14.48745,
  18.87931, 18.85293, 17.41729, 17.13374, 18.36859, 19.4126, 19.95924,
    20.37271, 21.50089, 19.26048, 15.43496, 15.92957, 16.62355, 17.5139,
    18.12078, 18.83948, 18.96633, 18.6112, 17.65306, 17.01452, 17.00873,
    16.78419, 16.73479, 16.36999, 16.09631, 17.47005, 17.78407, 16.26779,
    15.87397, 15.11122,
  19.0865, 19.90901, 19.54853, 19.12794, 19.39506, 19.80097, 20.67288,
    21.59486, 20.35263, 18.10597, 15.7552, 16.20699, 17.09133, 17.62681,
    17.74656, 18.38571, 18.42105, 18.21113, 17.93978, 17.15683, 17.05412,
    17.13203, 16.53424, 15.85085, 15.64049, 16.36259, 17.84193, 17.25902,
    16.03398, 15.21086,
  20.27496, 21.20519, 20.5433, 19.8097, 19.5083, 18.90774, 21.09083,
    22.31205, 19.04158, 16.35973, 16.12384, 16.77451, 17.36658, 17.46687,
    17.469, 17.7592, 17.83075, 17.85092, 17.76569, 17.00426, 17.00262,
    17.93449, 18.15186, 17.40201, 17.22834, 17.44175, 19.41622, 19.51446,
    16.24961, 14.55784,
  21.53877, 22.24971, 19.77969, 19.51397, 20.06133, 19.6042, 20.90926,
    20.55402, 16.80785, 15.65923, 16.11711, 16.72914, 16.94648, 17.0644,
    17.71364, 17.96673, 17.60772, 17.44779, 17.82292, 18.30429, 18.68711,
    18.9158, 18.69217, 18.17297, 18.12193, 18.35278, 19.01903, 20.8482,
    19.29748, 15.30289,
  20.39045, 19.33743, 19.18527, 21.42817, 22.31104, 22.12423, 21.44205,
    18.32241, 15.54727, 15.68256, 15.43337, 15.23128, 15.40277, 15.99101,
    17.22631, 18.11299, 18.35824, 18.77469, 18.7361, 18.4429, 18.59194,
    18.18418, 17.28077, 16.70954, 17.00624, 17.58466, 17.75392, 18.14598,
    18.72517, 16.25942,
  19.66989, 19.44691, 20.21058, 21.21593, 21.59208, 22.75307, 22.2082,
    18.06496, 15.27705, 15.7891, 15.91177, 16.26217, 16.8791, 17.574,
    18.37998, 19.27684, 19.12359, 18.27198, 17.75918, 17.06009, 16.5573,
    16.41574, 16.11641, 15.90022, 16.08182, 16.64968, 17.01154, 16.46199,
    15.88528, 14.8811,
  18.75929, 18.80801, 18.82804, 18.84921, 18.84236, 18.83092, 18.83719,
    18.85996, 18.86978, 18.89812, 19.63001, 19.96937, 18.98229, 19.14413,
    19.39642, 19.04618, 18.90756, 18.90817, 18.89623, 19.32944, 19.73735,
    19.31161, 19.20739, 19.62871, 19.75069, 19.3025, 21.48847, 24.14117,
    21.28034, 19.95924,
  19.02025, 19.16048, 18.90967, 19.20811, 19.05475, 18.83512, 18.87245,
    18.91199, 18.9679, 19.1308, 19.64044, 20.26849, 20.50379, 19.97809,
    19.60918, 19.75183, 19.07824, 19.00246, 19.38771, 19.96965, 20.0144,
    19.31931, 19.0238, 19.69426, 23.24375, 25.5641, 23.81377, 29.48981,
    23.15852, 20.95311,
  19.08596, 19.11093, 19.01234, 19.12542, 18.99806, 18.84469, 18.84632,
    18.93068, 19.04338, 19.1459, 19.26972, 19.75072, 20.22772, 20.56897,
    20.70313, 19.75553, 19.45565, 19.86457, 19.77977, 19.85859, 20.39568,
    21.55938, 22.44417, 21.81009, 26.9232, 33.81776, 27.66628, 29.7833,
    23.03063, 21.86705,
  19.05217, 18.99401, 19.15808, 19.31562, 19.47763, 19.93198, 19.95554,
    19.65828, 19.62317, 19.84953, 20.08272, 20.48578, 20.3846, 19.91001,
    20.93242, 21.79927, 21.34502, 19.99331, 19.57339, 19.42394, 21.75416,
    24.25248, 23.0027, 27.63074, 31.99809, 29.14716, 33.03787, 28.66471,
    22.91436, 20.87359,
  19.59424, 19.08298, 19.34417, 19.60005, 20.00692, 20.30986, 20.17504,
    19.8983, 20.46455, 21.51143, 21.74385, 21.13168, 20.26468, 20.51061,
    21.48534, 21.73483, 20.40572, 19.05166, 19.29784, 23.82176, 27.799,
    22.34602, 21.99584, 24.84875, 27.36197, 27.05353, 27.46266, 28.36656,
    28.3423, 22.19521,
  19.38636, 19.21736, 19.99368, 21.20398, 21.52822, 20.98457, 20.54991,
    20.3416, 20.14932, 20.37797, 20.28987, 21.5375, 23.91606, 24.04586,
    23.21058, 28.12603, 37.04298, 30.11109, 22.76735, 25.89145, 25.49249,
    20.77345, 21.47537, 22.52931, 25.13304, 25.8851, 26.13371, 40.71582,
    41.20353, 21.97857,
  19.24461, 19.56869, 20.59286, 21.97779, 22.57745, 21.96426, 21.56457,
    23.414, 23.87732, 23.61173, 24.22592, 24.42894, 23.49416, 22.9824,
    27.65183, 37.58701, 36.69099, 26.99689, 23.55395, 23.79865, 22.15482,
    20.85617, 21.50869, 24.01791, 26.27963, 23.70475, 30.03903, 51.48695,
    45.90335, 20.26136,
  19.34882, 19.81353, 20.92054, 22.19214, 22.09064, 23.57042, 26.33204,
    24.88935, 23.06737, 23.47586, 23.69168, 22.73477, 20.91579, 20.87387,
    24.34981, 28.41789, 25.83143, 23.72937, 22.11665, 21.91604, 21.42725,
    20.96688, 22.28318, 25.2847, 25.58918, 22.69683, 36.59001, 52.58826,
    30.17768, 20.30025,
  20.89632, 21.04811, 22.06135, 22.38525, 22.57561, 26.12832, 26.38309,
    22.95037, 22.95579, 23.47501, 22.81488, 21.26686, 20.32266, 23.89208,
    27.83088, 24.46872, 23.58154, 25.63091, 25.62463, 23.51868, 20.95875,
    22.18198, 26.5057, 28.68435, 24.36956, 24.17704, 33.58708, 37.26487,
    22.42834, 20.34414,
  22.74579, 23.36288, 25.91679, 29.45251, 29.19619, 26.60315, 22.11672,
    21.48627, 21.2244, 20.73645, 21.27353, 25.44704, 27.56614, 28.13227,
    27.26074, 26.93986, 27.92558, 28.86658, 27.98617, 26.0055, 25.77226,
    26.78247, 28.66768, 27.21736, 31.08676, 44.87746, 41.20878, 25.40187,
    21.12956, 19.27994,
  32.26848, 37.95948, 37.55751, 29.53958, 29.19935, 28.54945, 25.08493,
    26.24734, 28.16833, 32.40422, 39.28406, 29.03803, 25.98471, 25.5536,
    24.93785, 26.47787, 28.83826, 29.05805, 27.51154, 26.12672, 29.20622,
    29.80389, 26.55471, 23.306, 28.38302, 36.65045, 31.12488, 20.83538,
    19.76208, 18.87778,
  51.08892, 39.57608, 35.71294, 33.26972, 33.98859, 28.18068, 33.60141,
    34.30836, 28.77115, 33.40885, 35.78366, 23.20044, 24.34108, 26.19711,
    25.15429, 26.36015, 25.9685, 25.99635, 25.31919, 25.62006, 29.47939,
    28.92803, 23.09815, 26.11974, 31.79221, 25.40167, 20.38042, 19.86258,
    19.7543, 19.13305,
  65.08401, 49.22137, 52.91092, 60.19479, 62.87252, 58.14315, 49.21598,
    35.79651, 37.74342, 32.85783, 26.9501, 20.65308, 26.32854, 30.20933,
    27.16204, 25.63365, 26.31678, 25.50972, 24.43226, 27.73994, 31.14969,
    26.32817, 22.50676, 29.21277, 35.60506, 22.84021, 19.70429, 20.05394,
    20.37798, 19.6708,
  75.4543, 66.94144, 69.13499, 75.86205, 76.12899, 72.14072, 59.77184,
    55.64975, 46.30323, 35.06068, 41.73152, 42.69512, 48.10644, 49.91696,
    44.36295, 33.80801, 26.85801, 29.00937, 31.40243, 33.90737, 30.9844,
    26.92579, 31.88095, 29.39661, 25.52906, 20.67078, 19.76265, 19.69054,
    20.14113, 19.75384,
  51.09518, 63.16889, 78.55488, 84.08217, 82.42433, 70.75535, 69.49595,
    71.18198, 53.0055, 52.56016, 57.20009, 46.65894, 38.31654, 44.64666,
    48.71319, 33.08838, 31.56909, 32.25061, 34.61468, 37.1122, 33.43394,
    30.59695, 28.62667, 24.43967, 19.98105, 20.32775, 19.87503, 19.56055,
    19.5482, 19.31868,
  36.95411, 47.61491, 57.00178, 55.75051, 48.73298, 45.76284, 49.70552,
    41.31631, 38.41876, 41.9957, 42.10654, 32.63848, 27.25055, 33.51862,
    34.19272, 30.5585, 33.94098, 32.12552, 30.63182, 32.38472, 28.41784,
    25.68782, 22.43226, 21.26089, 20.72059, 20.34793, 19.89412, 19.67737,
    19.40857, 19.11482,
  30.56922, 31.77619, 31.4425, 28.61939, 26.12638, 28.47711, 30.59789,
    27.7528, 29.23237, 30.84502, 26.67251, 25.44807, 29.93502, 28.23122,
    29.18054, 30.75396, 32.52124, 29.71767, 29.06039, 31.32548, 23.41634,
    22.52489, 21.59455, 21.29391, 20.87387, 20.48071, 19.89887, 19.43708,
    19.25829, 19.0835,
  24.53678, 24.06911, 21.96028, 21.1847, 21.76497, 23.64444, 24.84969,
    25.4287, 25.64389, 23.75518, 22.444, 27.3857, 30.92027, 29.58111,
    35.5235, 34.7512, 30.34119, 26.02231, 28.87734, 30.18822, 22.391,
    22.3378, 21.57733, 21.51511, 20.49695, 20.15651, 19.93801, 19.17159,
    19.07811, 18.98388,
  23.62614, 22.99259, 20.52223, 19.68214, 20.37013, 21.03721, 21.82097,
    22.10777, 21.30836, 19.95819, 22.95903, 26.79806, 24.67153, 26.72009,
    31.76525, 30.85642, 29.59231, 28.20522, 31.1628, 30.70199, 25.00282,
    23.25021, 21.90983, 21.56072, 20.19426, 19.75462, 19.68157, 19.14867,
    19.02444, 18.9332,
  23.52601, 22.62133, 20.51335, 18.87023, 19.26964, 19.49611, 19.70481,
    19.63634, 19.04535, 21.29702, 25.30395, 23.42834, 21.35453, 23.05844,
    24.76063, 25.31635, 27.12438, 29.36649, 30.15246, 30.53412, 28.58132,
    26.02055, 22.33884, 21.59781, 20.54775, 19.77778, 19.53531, 19.20992,
    19.01297, 18.94461,
  22.37629, 22.01809, 20.19544, 18.6087, 18.6199, 18.81131, 18.71242,
    18.46788, 19.23612, 23.10526, 24.61333, 20.30602, 21.11072, 22.07648,
    22.26115, 22.74244, 24.03713, 25.49006, 26.02901, 26.97275, 28.24258,
    28.443, 24.1911, 22.43104, 21.04704, 20.18007, 19.56626, 19.2167,
    19.0222, 18.94786,
  23.40232, 21.49479, 19.98989, 18.94406, 18.93888, 18.22846, 18.27963,
    18.44934, 20.72062, 24.04329, 22.40725, 18.88588, 20.3279, 20.98496,
    21.16883, 21.82535, 22.50754, 22.86387, 23.72568, 24.24854, 26.15029,
    27.70514, 24.057, 24.66166, 23.17814, 21.00226, 19.70399, 19.35362,
    19.02818, 18.95312,
  23.51215, 21.77572, 19.93961, 18.67901, 19.39056, 19.63585, 19.84871,
    19.59919, 21.63662, 23.25183, 20.0059, 18.51581, 19.36566, 19.91723,
    20.13292, 21.45365, 22.59903, 22.34157, 22.52609, 22.57764, 24.34989,
    25.56497, 21.95638, 24.18215, 24.8348, 22.17378, 19.90624, 19.81429,
    19.35569, 18.9789,
  23.33871, 21.9091, 20.74505, 20.16349, 20.90443, 21.17484, 22.78055,
    24.17926, 25.49539, 22.843, 18.82919, 19.00679, 19.72775, 20.54527,
    20.89419, 22.05663, 23.43842, 23.20085, 22.34226, 22.51312, 23.5421,
    23.10666, 21.30071, 22.209, 23.42377, 23.49414, 21.76741, 20.2506,
    19.81182, 19.20516,
  22.73042, 22.8255, 20.86693, 20.17148, 21.71214, 23.36709, 24.10731,
    24.55339, 25.6964, 23.27002, 18.64016, 19.27752, 20.03474, 20.98677,
    21.62781, 22.84192, 23.61241, 23.77946, 22.99903, 22.3121, 22.41582,
    21.96976, 21.87288, 21.67144, 21.13043, 22.6036, 23.01299, 21.28354,
    20.73258, 19.95419,
  23.13757, 24.51133, 23.72361, 22.93536, 23.27274, 23.97005, 25.03303,
    26.13282, 24.41324, 22.08178, 19.12238, 19.74718, 20.69577, 21.18851,
    21.20205, 22.3692, 23.15278, 23.40943, 23.27249, 22.24502, 22.09099,
    22.27405, 21.67963, 20.79728, 20.42534, 21.2682, 22.94202, 22.46079,
    20.8818, 20.07462,
  24.68252, 26.15722, 25.07684, 23.56268, 23.28861, 22.9148, 25.73808,
    27.38382, 23.04519, 19.98624, 19.68187, 20.51817, 21.07499, 20.98458,
    20.90545, 21.7143, 22.5153, 22.97128, 23.06407, 22.03285, 22.06218,
    23.20208, 23.3695, 22.30235, 22.06832, 22.38755, 24.58074, 24.9323,
    21.16419, 19.27971,
  26.88663, 29.12529, 23.73153, 22.86364, 23.75453, 23.56707, 25.29507,
    25.11633, 20.47928, 19.14876, 19.82302, 20.51913, 20.59112, 20.52061,
    21.22108, 21.94366, 22.19581, 22.46805, 23.00171, 23.34186, 24.00857,
    24.57895, 24.04775, 23.26129, 23.01316, 23.39798, 24.2906, 26.25973,
    24.59224, 20.15186,
  24.90906, 23.64967, 22.80791, 26.97671, 27.73208, 26.4756, 26.08924,
    22.39273, 19.03079, 19.21249, 19.06758, 18.78159, 18.79976, 19.23805,
    20.54557, 21.92119, 22.85223, 23.87873, 24.03651, 23.61614, 23.97025,
    23.66253, 22.4478, 21.67311, 21.91719, 22.6109, 22.9124, 23.38128,
    23.90576, 21.28196,
  23.26144, 22.86562, 24.74917, 27.52164, 27.52925, 28.01246, 27.17693,
    22.24439, 18.80368, 19.44097, 19.60915, 19.90405, 20.39347, 20.88744,
    21.73661, 23.15672, 23.69185, 23.38821, 22.98228, 22.14768, 21.61109,
    21.41366, 21.00391, 20.70607, 20.93155, 21.59097, 21.99906, 21.44607,
    20.82319, 19.67256,
  27.02094, 27.10463, 27.17191, 27.23054, 27.20054, 27.20708, 27.2552,
    27.31155, 27.37053, 27.64832, 29.0656, 29.74203, 27.66157, 28.00703,
    28.42944, 27.67181, 27.38626, 27.43493, 27.56657, 28.18906, 28.69143,
    28.48982, 28.9708, 29.85274, 30.51724, 30.92393, 34.72855, 39.00788,
    32.27848, 29.53853,
  27.60293, 27.92519, 27.38483, 27.90987, 27.61753, 27.27029, 27.41174,
    27.56666, 27.76714, 28.15676, 29.06485, 30.18696, 30.7114, 29.63919,
    28.74873, 29.07757, 27.78355, 27.84333, 28.74585, 29.75324, 29.63691,
    28.93251, 29.31106, 32.25024, 39.67628, 45.15569, 40.47884, 47.94527,
    35.25961, 31.00336,
  27.5822, 27.63762, 27.5076, 27.62034, 27.45059, 27.31849, 27.39299,
    27.6117, 27.81814, 27.98552, 28.28828, 29.12278, 29.92036, 30.61193,
    30.93975, 29.16634, 28.78178, 29.61347, 29.59056, 30.19297, 32.16217,
    35.80996, 38.1111, 39.06099, 48.78205, 58.34878, 49.15595, 48.65308,
    35.38425, 32.72717,
  27.55015, 27.56954, 27.96582, 28.37338, 28.65045, 29.45648, 29.56993,
    29.0641, 29.05489, 29.63203, 30.16164, 30.74047, 30.50594, 29.65019,
    31.67967, 33.45646, 32.53215, 30.00216, 30.12931, 31.64202, 37.09026,
    41.722, 40.99165, 49.64425, 55.0106, 49.83503, 57.49546, 46.09697,
    35.45869, 30.75459,
  28.53443, 27.86214, 28.58467, 29.28785, 29.95501, 30.06557, 29.70406,
    29.6225, 31.1216, 32.78127, 31.98536, 31.0361, 30.2549, 31.14171,
    32.54607, 33.23418, 32.27785, 30.00137, 32.07632, 39.79784, 45.54183,
    37.24602, 38.07576, 41.79172, 43.03718, 43.74443, 44.90383, 49.5136,
    45.86359, 31.98616,
  27.99516, 28.44366, 30.22946, 32.31088, 32.05416, 30.61204, 30.31947,
    29.98676, 29.54803, 29.94736, 30.09918, 33.1795, 38.13274, 38.50326,
    41.47217, 49.32869, 56.15977, 48.98985, 39.93179, 43.24881, 40.53262,
    33.76602, 35.29844, 37.64966, 41.02878, 42.37769, 47.25518, 69.06816,
    62.84155, 31.15788,
  27.60584, 28.75756, 30.81583, 32.96461, 32.98334, 31.90204, 33.19011,
    37.35502, 38.25399, 36.95932, 37.64766, 37.83506, 35.82016, 37.47939,
    45.4945, 55.42806, 51.99466, 43.48724, 38.64681, 38.30639, 35.15149,
    33.45803, 35.30503, 40.49411, 45.31216, 43.26685, 53.3228, 76.70195,
    63.24084, 29.11869,
  26.82697, 28.19025, 30.53401, 32.8246, 32.88903, 36.48916, 42.01557,
    38.32604, 34.61081, 34.97921, 34.39452, 32.44136, 30.1586, 32.19679,
    37.11125, 41.37867, 39.86263, 38.56686, 34.81401, 34.45555, 33.41355,
    33.08808, 36.5435, 42.31941, 43.18626, 40.67448, 55.47853, 70.47787,
    41.44552, 29.93984,
  28.07589, 28.57611, 31.174, 32.7606, 34.2098, 39.15788, 37.41993, 32.83539,
    33.22821, 33.09221, 31.08599, 29.01782, 28.91483, 36.31815, 44.12995,
    38.3718, 37.28939, 41.48369, 42.0651, 37.90798, 33.29699, 37.35979,
    46.51226, 49.72312, 41.45337, 43.1053, 51.98098, 55.59743, 33.62038,
    29.62331,
  32.46189, 35.98031, 38.76475, 44.44133, 43.70005, 38.92506, 27.85151,
    27.56104, 26.57725, 27.26737, 30.48383, 39.12341, 43.1289, 43.45068,
    41.60942, 41.9723, 44.98508, 48.01966, 43.42761, 39.26107, 40.24704,
    42.1627, 44.8499, 45.16148, 55.17054, 71.21626, 60.36008, 37.64962,
    30.08778, 27.55143,
  51.05629, 53.83961, 53.11821, 45.9998, 44.13423, 40.65448, 34.33857,
    38.04497, 43.65665, 50.30906, 58.42198, 42.12321, 36.18867, 35.9892,
    36.6406, 40.1013, 44.27322, 44.38941, 41.42099, 40.00973, 43.12423,
    44.07864, 39.25679, 37.01654, 44.23048, 50.14498, 41.17361, 29.03595,
    28.22985, 27.09661,
  72.48426, 53.61577, 53.85674, 54.67653, 55.3855, 46.25026, 53.72002,
    54.31546, 48.40612, 50.25832, 46.64284, 32.39956, 34.66436, 37.45417,
    37.14798, 39.943, 39.87206, 39.80244, 39.05395, 40.85703, 44.34304,
    41.59238, 34.55003, 39.63124, 45.98207, 35.64103, 28.79278, 28.51924,
    28.37523, 27.50073,
  87.55037, 76.05486, 92.17421, 101.6797, 102.5294, 90.28004, 72.39165,
    54.05697, 55.86363, 43.76408, 36.58237, 32.71471, 41.04041, 46.44514,
    43.3377, 39.5928, 40.36691, 39.62856, 38.66163, 45.93752, 49.26958,
    37.92292, 34.70849, 41.54308, 46.51185, 31.77189, 28.17171, 28.90844,
    29.22326, 28.27395,
  107.3475, 119.0432, 118.7079, 117.3578, 105.6889, 95.75096, 85.84797,
    80.80563, 63.59245, 55.41747, 68.93768, 68.09573, 73.95203, 76.44478,
    66.59329, 50.28258, 43.19927, 46.83534, 51.5715, 54.13865, 47.76846,
    40.60612, 45.9537, 39.56571, 33.36129, 29.49385, 28.49016, 28.26443,
    28.74986, 28.29241,
  88.91507, 89.41611, 88.56315, 84.62068, 76.49535, 77.69511, 97.48117,
    95.28802, 79.5061, 85.03845, 87.35715, 73.66251, 67.67048, 73.38216,
    71.35854, 55.40355, 53.03227, 56.22857, 61.24835, 62.00792, 50.70922,
    46.46982, 40.40401, 33.18011, 28.72886, 29.25, 28.55028, 28.04312,
    27.9417, 27.65299,
  74.44976, 71.48287, 70.63698, 66.90977, 72.15856, 82.10054, 82.10799,
    77.26894, 70.97135, 72.49756, 68.97412, 58.58532, 52.5427, 59.58939,
    57.38676, 54.73286, 57.68243, 55.79567, 56.46969, 56.5768, 42.03225,
    36.8187, 32.27257, 30.57369, 29.94683, 29.28267, 28.50681, 28.16398,
    27.8143, 27.43501,
  59.07769, 55.7011, 52.14098, 54.60313, 57.75247, 57.96008, 61.26826,
    67.32314, 57.01648, 55.45398, 50.16951, 48.47358, 53.99023, 51.85524,
    53.63919, 53.87333, 54.26316, 50.31292, 51.76269, 51.75511, 33.97112,
    31.42855, 31.05929, 31.45325, 30.19534, 29.35716, 28.52116, 27.81937,
    27.60358, 27.39677,
  43.24741, 41.81735, 39.50218, 42.06676, 45.15286, 49.96323, 55.10947,
    54.16032, 46.04776, 41.82431, 44.03626, 54.8469, 58.70369, 58.9439,
    63.80719, 57.93021, 48.73029, 43.46744, 49.17499, 47.1167, 32.28035,
    33.09791, 32.58212, 31.93999, 29.29695, 28.84328, 28.55582, 27.47805,
    27.35531, 27.2539,
  39.01877, 38.39671, 35.25546, 34.93159, 38.50028, 43.0265, 43.72277,
    39.73526, 35.68157, 35.66208, 44.67445, 53.35434, 50.46378, 54.98185,
    56.57878, 48.39078, 46.53533, 49.24007, 54.17664, 49.53988, 38.22292,
    36.51469, 33.75329, 31.72085, 28.77044, 28.40533, 28.23494, 27.48197,
    27.30174, 27.20028,
  38.85143, 37.87566, 34.52644, 31.78584, 34.0967, 35.16336, 33.66786,
    31.45665, 31.61872, 39.41663, 48.30848, 45.10906, 43.85159, 45.94758,
    43.43954, 39.67554, 42.34847, 49.32248, 52.23091, 51.46828, 46.84599,
    41.13609, 34.25294, 31.78095, 29.46483, 28.53022, 28.07973, 27.60856,
    27.33059, 27.23788,
  36.99509, 37.16443, 32.63868, 29.69103, 30.80437, 30.76079, 29.17887,
    29.08669, 32.73929, 41.76125, 44.42917, 38.31488, 41.24416, 39.37607,
    36.43972, 35.81238, 38.66684, 43.29876, 45.12228, 46.03801, 45.70222,
    43.63203, 36.86075, 32.99927, 29.99592, 29.01842, 28.10495, 27.63668,
    27.37195, 27.27131,
  38.21489, 35.22342, 31.54407, 29.53737, 29.73901, 27.69815, 28.01131,
    29.52074, 35.54253, 42.4593, 39.63203, 34.5129, 36.2516, 33.74632,
    32.19549, 33.22434, 35.5409, 38.09622, 40.05951, 41.15342, 42.21873,
    42.20254, 38.47171, 37.50449, 34.08315, 30.42436, 28.35732, 27.8663,
    27.39921, 27.27089,
  37.29203, 34.72504, 30.54845, 27.92508, 29.63297, 30.31953, 31.39625,
    31.67882, 36.66749, 40.51061, 34.2779, 30.84241, 30.74952, 30.13709,
    29.58852, 32.05838, 34.99765, 35.51025, 36.99925, 38.30983, 38.97898,
    38.80179, 36.0129, 37.88351, 37.5741, 32.57374, 28.73453, 28.68561,
    27.89566, 27.34154,
  37.33375, 34.76749, 32.47451, 31.39813, 32.93246, 33.6725, 37.19004,
    38.27152, 41.5596, 38.98591, 30.58892, 29.6808, 30.5478, 31.58203,
    31.58813, 33.80011, 36.47899, 36.71213, 36.78825, 37.46976, 36.69551,
    35.4044, 34.68095, 35.92184, 36.72519, 35.59739, 32.05099, 29.34409,
    28.47156, 27.63647,
  35.19358, 37.18887, 31.70044, 30.87723, 34.33072, 36.96056, 38.41403,
    39.03151, 42.46854, 38.5579, 28.85016, 29.5155, 30.95643, 32.91437,
    33.8627, 36.05108, 36.92289, 37.4991, 36.66628, 34.39999, 34.663,
    35.49793, 35.01231, 33.54575, 32.01192, 33.53896, 33.50396, 30.69191,
    29.81412, 28.74042,
  37.20357, 41.37537, 38.22254, 36.51008, 37.49574, 38.00657, 39.37226,
    41.31545, 40.67863, 35.87958, 29.32211, 30.66388, 32.87017, 34.00864,
    33.83094, 35.62835, 36.26962, 36.6053, 35.62635, 32.96636, 34.78123,
    36.55073, 33.67841, 30.7118, 29.68534, 31.06891, 33.09369, 32.34694,
    29.99398, 28.85684,
  41.60061, 45.92943, 42.17157, 38.07201, 39.17854, 38.0642, 40.93106,
    42.05964, 36.68449, 31.39124, 30.69935, 32.62635, 34.18386, 33.88086,
    33.60409, 34.40714, 35.07118, 35.43667, 34.72009, 32.55014, 34.66386,
    37.49527, 35.84107, 32.9121, 31.95182, 32.82895, 35.66473, 35.90454,
    30.37926, 27.71367,
  46.38663, 49.75278, 40.56721, 37.81086, 41.34263, 40.21227, 42.30019,
    40.42371, 31.24645, 30.25372, 32.11019, 33.1162, 33.60598, 33.86762,
    34.64244, 34.4842, 33.91969, 34.23746, 34.43753, 34.46086, 37.89639,
    40.25169, 36.95457, 34.41226, 33.3094, 34.23876, 35.50067, 37.94208,
    35.28757, 28.95858,
  40.05966, 34.35915, 34.93976, 42.90269, 44.51756, 44.72404, 44.10614,
    35.87156, 28.79903, 30.44567, 30.39725, 29.60538, 30.3283, 31.98765,
    33.73833, 34.28342, 34.99692, 37.1148, 36.63199, 35.04553, 36.83633,
    36.41257, 33.39293, 31.69733, 31.86236, 32.97354, 33.47169, 33.96331,
    34.11308, 30.57746,
  35.94662, 34.79943, 39.59752, 43.37915, 42.34364, 45.1052, 46.671,
    35.62886, 28.8554, 30.9614, 31.49994, 33.15001, 34.87329, 35.65083,
    36.23144, 37.01104, 37.08959, 36.24467, 34.76878, 32.6643, 32.0266,
    31.18857, 30.47119, 30.05285, 30.43311, 31.31049, 31.78773, 30.99296,
    29.85972, 28.2057,
  31.08328, 31.57352, 32.10054, 32.69781, 33.05574, 33.54901, 34.15342,
    34.82081, 35.66176, 37.20391, 40.01368, 40.41308, 35.74153, 37.0609,
    37.82201, 36.86073, 37.85327, 40.11906, 42.97609, 47.1336, 49.97702,
    49.44122, 51.50317, 55.25499, 58.19388, 58.75069, 63.76482, 65.27403,
    42.31888, 35.62332,
  32.53008, 33.21815, 32.2173, 33.7035, 33.22823, 33.24854, 34.2503,
    35.12982, 36.19163, 37.68293, 40.00103, 43.11821, 44.94444, 42.46041,
    41.4748, 43.79535, 43.06014, 46.42328, 50.66984, 54.45399, 55.75785,
    56.61476, 59.7742, 67.61156, 74.73085, 69.73791, 62.72915, 66.37611,
    44.22331, 37.74667,
  30.22457, 30.47915, 30.95954, 31.47602, 31.91405, 32.60762, 33.38328,
    34.39038, 35.58206, 36.9981, 38.97536, 42.21797, 45.95972, 50.27048,
    53.63132, 52.6261, 56.06625, 60.98949, 65.05911, 71.36443, 79.9286,
    87.97853, 91.23714, 92.23814, 91.87885, 83.41101, 76.8643, 64.13631,
    44.88547, 40.02796,
  33.71346, 34.75421, 36.74805, 38.83637, 40.6523, 42.88802, 43.30254,
    42.96851, 44.24222, 46.41465, 48.02084, 50.07578, 52.15327, 54.1045,
    61.81087, 66.60813, 65.0661, 63.60375, 70.51231, 78.69443, 89.41331,
    92.1768, 89.09982, 96.22865, 94.78699, 92.46268, 82.81389, 63.50606,
    45.03106, 36.57357,
  37.96972, 37.04563, 39.60636, 41.30609, 42.87381, 43.26768, 43.85761,
    45.41508, 48.96075, 52.17385, 52.49432, 54.57411, 57.08049, 61.064,
    65.03978, 67.60257, 66.70285, 63.55582, 69.33073, 79.59782, 82.53546,
    73.44539, 75.26037, 84.44273, 90.79713, 89.77244, 83.64061, 88.97814,
    75.16617, 44.77284,
  39.42572, 42.50874, 46.96346, 51.91979, 52.14356, 51.32307, 54.77838,
    57.85629, 60.7084, 66.3046, 74.5133, 87.1722, 100.0688, 99.9863,
    105.3643, 112.086, 107.0651, 93.96893, 81.18054, 80.67183, 74.3493,
    66.55273, 73.99812, 81.62306, 89.94342, 91.12996, 89.72478, 103.5026,
    85.71046, 42.5996,
  46.01919, 52.32457, 59.16663, 66.86079, 71.60242, 76.53369, 84.93966,
    94.04225, 94.56564, 91.59372, 89.34224, 83.21274, 74.3499, 76.83406,
    80.90836, 85.20747, 86.05457, 77.37143, 66.44012, 69.26859, 67.13004,
    67.73219, 74.65523, 84.13036, 86.41704, 78.8569, 84.56736, 93.2815,
    70.55505, 34.75964,
  52.89593, 59.9409, 67.145, 74.22667, 76.63857, 83.96348, 88.03561,
    70.41254, 59.45118, 59.35928, 55.72416, 52.46264, 49.64525, 52.69243,
    57.35002, 63.95, 67.70087, 67.33031, 61.50376, 63.61047, 64.51794,
    68.39938, 76.9599, 83.53473, 79.9348, 76.84859, 87.87363, 84.74611,
    58.85292, 35.71692,
  63.17144, 65.71138, 69.97977, 71.68071, 69.67358, 72.48253, 63.778,
    59.99038, 63.0373, 64.77241, 65.5246, 66.51011, 71.33668, 85.86807,
    95.02405, 78.5941, 80.41298, 87.66586, 88.35047, 81.05762, 78.15388,
    91.70743, 104.8407, 103.6373, 88.57471, 94.65722, 92.57957, 75.15402,
    42.7487, 35.45942,
  88.28866, 95.1306, 91.81998, 95.43392, 86.66957, 75.9274, 60.67982,
    70.94006, 74.83966, 86.54606, 99.93346, 112.8032, 110.8785, 106.2653,
    100.2722, 108.7623, 112.6023, 110.8577, 104.8746, 102.3877, 109.5784,
    106.2426, 100.2884, 89.89656, 95.21124, 103.9724, 85.59155, 51.48993,
    35.18237, 32.04248,
  113.1068, 106.662, 108.2177, 98.68056, 110.5999, 111.9728, 108.3757,
    112.8558, 117.8319, 119.4146, 109.817, 83.84729, 82.60316, 84.47451,
    88.98625, 95.09969, 100.1288, 99.12088, 95.67446, 95.36237, 104.8219,
    97.71137, 75.02089, 67.43766, 74.02542, 71.62879, 50.83252, 35.35657,
    34.31632, 31.89398,
  124.6622, 108.8077, 120.2554, 125.6304, 117.9881, 100.5538, 101.6121,
    94.48812, 85.10921, 75.20373, 70.02177, 68.15317, 76.04406, 83.36786,
    85.4965, 84.89336, 82.16161, 81.27379, 78.66976, 80.56951, 89.87821,
    82.24585, 63.4234, 73.05341, 74.67647, 54.13713, 35.2251, 37.72992,
    35.48935, 33.22991,
  147.6759, 148.4615, 150.9646, 150.7524, 148.9241, 127.6895, 103.829,
    96.35127, 97.57822, 77.04558, 77.02531, 78.70576, 91.45491, 101.0779,
    94.86292, 80.08235, 82.3562, 79.49155, 77.91191, 85.25075, 88.08919,
    75.20767, 67.24217, 64.90024, 60.57929, 46.68066, 37.1254, 39.16185,
    38.09254, 35.08774,
  145.7521, 145.9906, 145.1566, 140.8969, 132.1719, 137.9812, 142.8965,
    143.8526, 126.931, 131.9564, 143.4789, 137.1772, 144.9353, 147.8364,
    125.4552, 104.5164, 102.8146, 108.2198, 112.679, 106.3575, 88.1696,
    68.98272, 62.93672, 50.83406, 43.35317, 40.5154, 37.11024, 36.02483,
    35.87554, 34.45022,
  106.6809, 101.8306, 106.5294, 111.5831, 119.813, 135.0318, 147.3672,
    148.9433, 146.0765, 147.0239, 143.5932, 136.3942, 142.2929, 145.2513,
    139.6395, 134.9683, 120.2621, 115.6356, 112.3771, 99.88084, 65.89212,
    60.47527, 49.04188, 42.52292, 40.21099, 38.50895, 36.23178, 34.61855,
    33.68317, 32.86596,
  100.4715, 106.3192, 111.8154, 116.237, 119.8418, 129.459, 140.7745,
    132.3259, 124.1975, 123.5499, 124.5897, 118.156, 116.343, 130.2867,
    125.6875, 118.3325, 113.3106, 96.40562, 85.90225, 73.57741, 50.4071,
    49.91838, 43.15913, 41.75291, 40.24601, 37.95599, 35.64036, 34.72518,
    33.5032, 32.62317,
  90.81255, 89.3745, 92.16626, 95.74105, 99.61047, 104.4338, 109.1327,
    110.9391, 109.3633, 109.1611, 105.1992, 117.9032, 132.6624, 121.4855,
    113.271, 104.0485, 93.20141, 79.68809, 75.42802, 69.14108, 46.5028,
    48.32367, 44.08587, 42.03274, 39.78162, 38.29999, 35.46603, 33.48809,
    32.92394, 32.51325,
  72.69556, 75.91603, 75.72601, 80.215, 84.79264, 91.13451, 95.86486,
    99.61814, 103.6989, 106.6504, 122.24, 142.0402, 140.8276, 133.3485,
    126.522, 101.7708, 79.20837, 69.62228, 75.54674, 68.90843, 48.72962,
    49.62077, 45.00988, 42.89355, 38.4725, 36.69331, 35.29064, 32.57018,
    32.3542, 32.11833,
  80.37897, 76.48113, 67.14191, 64.83993, 70.35641, 75.46004, 82.32505,
    90.34856, 96.04933, 105.6093, 120.331, 120.3054, 102.6427, 103.0146,
    97.69511, 90.69353, 92.15302, 95.59409, 95.07346, 81.48523, 59.15869,
    51.62773, 45.7092, 41.73623, 37.14601, 35.46688, 34.44595, 32.70962,
    32.24273, 32.09254,
  75.92094, 68.99092, 59.47467, 54.42271, 60.59208, 67.07249, 75.06573,
    82.84399, 91.37699, 102.5875, 104.5158, 85.63737, 80.38766, 81.06772,
    80.36031, 81.93123, 88.90622, 95.51779, 93.30912, 85.81687, 71.33216,
    57.99039, 46.68366, 42.40925, 38.96552, 35.92158, 34.46806, 32.99899,
    32.22683, 32.14153,
  67.60646, 60.93, 52.80339, 50.62796, 56.64106, 63.36994, 69.45039,
    75.29362, 81.88461, 88.15266, 80.81137, 66.87804, 75.64684, 77.54837,
    77.39589, 76.78947, 78.19159, 78.15132, 76.97585, 73.29974, 68.13445,
    64.05342, 54.54465, 46.94021, 41.39892, 37.45923, 34.52306, 33.07019,
    32.28713, 32.17578,
  68.67236, 58.22134, 53.84337, 53.11802, 58.68361, 59.99651, 65.5649,
    68.64596, 75.987, 78.48313, 67.10757, 62.61896, 71.47167, 72.74522,
    71.26407, 69.36244, 66.37814, 63.82111, 63.36332, 62.23346, 61.43994,
    60.3301, 58.21659, 56.15556, 48.20556, 38.98776, 34.70677, 33.5539,
    32.37548, 32.17007,
  66.86473, 61.49032, 54.63253, 54.93276, 64.2809, 68.10443, 68.44022,
    65.32779, 67.84106, 65.90931, 55.14189, 59.24733, 64.58238, 65.94939,
    63.71248, 62.79868, 60.71202, 56.12496, 54.82399, 54.94632, 55.09164,
    54.58625, 52.79378, 53.49773, 52.25996, 42.89168, 36.59261, 35.95312,
    33.78298, 32.31415,
  74.59705, 71.68108, 70.05071, 72.76016, 77.2795, 76.53384, 78.27982,
    75.44177, 75.52029, 65.6424, 54.70916, 63.68547, 68.01521, 70.31233,
    67.45379, 65.26068, 63.48689, 58.65662, 54.26035, 53.46305, 53.03763,
    51.54208, 50.08435, 49.66278, 50.49017, 49.60494, 43.45488, 37.28457,
    35.34416, 33.13284,
  77.63773, 81.58257, 73.42802, 74.79765, 78.20792, 77.77148, 74.51272,
    74.59296, 79.54719, 70.75565, 57.61861, 66.78876, 70.07635, 72.14077,
    70.11359, 68.43349, 64.02641, 60.30435, 56.1111, 52.60522, 52.59389,
    52.63259, 49.98956, 47.19153, 46.28699, 49.16221, 49.04716, 42.6218,
    39.24202, 35.97586,
  91.68073, 97.2958, 92.70847, 85.81441, 81.0376, 76.79329, 81.31831,
    85.70938, 79.73245, 68.53619, 66.68231, 72.37569, 74.78534, 72.91219,
    67.82216, 65.73206, 63.16642, 60.4044, 57.91151, 54.05515, 53.5342,
    52.35936, 47.85317, 44.85592, 45.60451, 48.28444, 51.0549, 46.99006,
    38.81612, 35.52073,
  103.2638, 102.9513, 91.54821, 82.20411, 78.6728, 76.37551, 84.61818,
    84.80255, 71.3807, 66.61021, 72.46455, 75.93262, 74.97464, 70.9455,
    66.99602, 63.5859, 60.61659, 57.95045, 55.95205, 53.36609, 55.29108,
    58.81879, 58.0774, 54.81241, 54.42904, 56.25725, 59.14396, 54.31813,
    39.69958, 33.06009,
  104.4236, 98.95156, 88.25726, 88.27238, 88.64492, 85.00134, 86.29419,
    78.58717, 65.69939, 69.79563, 74.19297, 74.83032, 73.10223, 69.71518,
    67.13389, 63.19127, 58.67388, 58.07244, 60.91454, 64.37698, 66.94744,
    66.08781, 61.29931, 58.80573, 58.60286, 60.08652, 60.67359, 61.64787,
    52.93883, 36.67496,
  84.11077, 81.88705, 91.05109, 98.24259, 97.64955, 96.26271, 87.66969,
    67.31815, 61.36913, 64.34496, 61.96067, 61.07555, 62.17092, 63.98216,
    66.47781, 67.5005, 68.00858, 69.815, 68.57056, 65.25047, 63.86848,
    60.05583, 55.40586, 52.95847, 53.59773, 54.37066, 53.41824, 50.48893,
    47.69466, 40.16584,
  87.41539, 90.93336, 91.47142, 90.3229, 91.04539, 96.35761, 91.36356,
    69.44632, 59.7461, 65.7427, 69.94978, 75.37018, 78.72527, 79.04781,
    76.50388, 74.51828, 68.19177, 61.66983, 58.28071, 54.71317, 51.43218,
    49.40512, 47.67378, 46.48349, 46.21436, 46.31891, 45.01675, 41.03051,
    37.17044, 33.0533,
  38.05968, 39.2006, 40.37812, 41.85604, 43.20258, 44.83866, 46.64091,
    48.52912, 50.55983, 53.01573, 56.33143, 57.6069, 54.84675, 55.85497,
    56.4233, 55.48223, 55.02763, 55.19404, 55.48057, 56.58239, 56.85792,
    55.12461, 55.76598, 58.0903, 59.11926, 57.41383, 60.03278, 61.45052,
    45.84362, 40.79541,
  41.80123, 43.83454, 44.61344, 47.20733, 48.41796, 50.07, 52.42911,
    54.85724, 57.40495, 60.13742, 63.33628, 66.92974, 69.12193, 67.73075,
    66.95435, 67.72392, 66.29245, 67.27182, 68.77785, 70.23598, 70.04584,
    68.96314, 68.58265, 70.91823, 73.35175, 66.5364, 57.10155, 59.92839,
    46.57393, 42.23317,
  45.35759, 47.82641, 49.91343, 51.97639, 53.65559, 55.26128, 56.72771,
    58.34168, 60.14222, 61.86524, 63.65138, 66.02221, 68.20021, 70.58455,
    72.00929, 69.71913, 70.64477, 73.0779, 75.56757, 80.05074, 86.65759,
    92.15156, 92.12788, 88.60287, 84.50539, 78.35825, 69.89663, 58.14391,
    45.73383, 42.91483,
  52.62685, 55.47293, 58.54609, 61.54762, 64.03189, 66.41528, 67.19903,
    67.38342, 68.56688, 69.55371, 69.90311, 70.59517, 70.16658, 69.16472,
    72.21046, 73.65607, 70.11568, 67.76074, 72.19747, 77.40176, 85.21455,
    86.79899, 83.58366, 88.75616, 87.25907, 85.51755, 81.07348, 65.62846,
    50.58769, 41.89827,
  63.166, 64.76762, 67.936, 70.31609, 71.87527, 72.89954, 74.07394, 74.86938,
    77.02246, 78.80803, 79.20951, 82.25209, 83.85641, 83.06087, 82.60652,
    81.92946, 77.6482, 71.65913, 72.21474, 77.19455, 76.76464, 68.36932,
    70.5383, 77.32188, 83.42097, 85.0524, 82.12675, 87.61813, 77.37752,
    50.02877,
  71.35274, 75.72813, 79.61227, 83.4295, 82.84651, 81.82233, 84.57585,
    84.82478, 83.47902, 84.44223, 88.49954, 97.60706, 107.0359, 104.3548,
    104.0471, 104.9746, 102.4234, 92.80437, 81.44979, 78.65358, 70.68135,
    63.08748, 68.0894, 72.34778, 76.62277, 76.51798, 76.43668, 89.26061,
    80.76561, 46.03713,
  68.3688, 73.00286, 77.60509, 82.41225, 84.58958, 87.67665, 94.29551,
    99.29699, 97.98427, 92.80319, 88.64088, 80.62455, 71.83047, 74.26677,
    76.26547, 78.86903, 79.53287, 75.89063, 70.26633, 71.05975, 68.71791,
    67.94164, 71.39275, 76.41638, 76.21262, 70.32092, 72.968, 79.09722,
    66.90393, 39.50348,
  66.92998, 72.407, 78.45793, 84.20426, 87.53102, 95.66006, 99.87513,
    85.52722, 79.20802, 81.98883, 81.08018, 79.75183, 78.86032, 79.911,
    80.10902, 80.79192, 82.07465, 79.79932, 74.34718, 73.54981, 74.06107,
    77.03547, 81.39514, 82.39909, 77.10693, 75.05106, 81.01108, 77.10951,
    56.98993, 40.92229,
  87.3951, 91.06298, 94.45043, 97.50325, 98.97676, 102.1194, 95.18953,
    96.25443, 100.5856, 103.5502, 104.9362, 104.7945, 105.6631, 111.8297,
    113.3927, 99.6143, 96.98134, 97.62236, 94.04464, 85.86766, 81.95245,
    88.39944, 95.46626, 92.29364, 81.7705, 85.27547, 82.4361, 67.26074,
    43.22522, 40.39438,
  120.1619, 125.0613, 117.573, 117.5013, 117.1031, 110.0234, 92.23961,
    98.48444, 96.97816, 99.75195, 103.581, 108.7557, 105.5948, 99.64168,
    94.80946, 99.52449, 101.0799, 99.13186, 95.08919, 93.51189, 94.81168,
    88.91972, 82.09541, 73.91562, 77.62592, 84.68831, 73.45822, 50.22161,
    39.93402, 38.07281,
  145.1018, 140.4838, 136.9249, 123.4136, 127.477, 119.6023, 109.44,
    108.3187, 106.8096, 100.7052, 87.13539, 70.32491, 68.01205, 68.31773,
    68.84033, 70.58128, 73.73935, 75.22426, 76.00169, 80.02229, 89.01366,
    82.77142, 68.28958, 65.57057, 69.48898, 65.74001, 50.24141, 40.92902,
    40.33361, 38.27945,
  152.6227, 147.8153, 149.5591, 148.6593, 143.8123, 118.8317, 111.6687,
    102.1481, 93.13116, 84.21205, 79.11177, 75.37031, 77.48499, 77.5959,
    73.09949, 70.00536, 67.95729, 68.11671, 68.80223, 72.80478, 80.70778,
    77.71077, 66.07025, 74.12093, 75.62384, 59.71547, 42.18818, 45.7294,
    42.00773, 39.6993,
  155.5734, 155.4317, 156.6446, 156.8486, 155.1258, 150.0906, 141.0435,
    127.3286, 131.8684, 115.0404, 109.2687, 101.4833, 106.6125, 107.0133,
    93.19574, 76.45297, 76.82198, 74.78127, 73.23936, 76.58086, 76.99874,
    69.05545, 61.96245, 57.08094, 56.17183, 51.17539, 42.92069, 44.32748,
    43.84496, 41.05489,
  142.3198, 143.6363, 142.5671, 143.4554, 143.0531, 143.1913, 143.5576,
    142.5944, 138.8053, 137.8938, 137.2656, 134.385, 135.1045, 135.1729,
    118.2814, 94.51385, 87.47156, 89.56258, 90.68868, 82.72124, 70.01663,
    60.94836, 55.05694, 47.1368, 43.27457, 43.05921, 41.28169, 40.32484,
    40.78061, 40.10006,
  111.9134, 110.8914, 115.4684, 119.0634, 121.3082, 123.1504, 127.8902,
    123.1678, 114.9169, 112.7522, 106.254, 100.6221, 103.6152, 106.2127,
    103.578, 100.2488, 88.24792, 82.3168, 80.93736, 74.58902, 56.88231,
    56.06524, 49.1029, 46.00251, 44.85461, 43.13938, 41.66075, 40.41536,
    39.34324, 38.7839,
  111.3343, 115.9378, 116.8962, 116.1857, 113.6072, 113.9079, 114.3423,
    105.881, 95.02662, 89.51692, 88.25831, 83.73983, 80.63754, 88.01051,
    85.32911, 82.63466, 81.77724, 72.99764, 69.2774, 62.89822, 50.57829,
    51.75346, 47.4689, 46.04901, 44.97883, 43.19562, 41.21377, 40.53689,
    39.52647, 38.76539,
  95.88968, 95.27622, 97.29668, 99.56396, 100.7625, 102.0871, 103.2966,
    102.2506, 98.56234, 93.47569, 87.6051, 95.08205, 101.227, 92.9422,
    86.17896, 80.22287, 73.45532, 68.49955, 68.23279, 62.8424, 50.02848,
    51.49741, 47.98671, 45.71262, 44.2617, 43.18593, 40.65709, 38.97025,
    38.81057, 38.5725,
  88.98273, 91.03662, 89.02496, 90.61768, 91.9633, 94.07887, 94.4169,
    95.11713, 97.06352, 98.22997, 108.0943, 116.0893, 112.3575, 107.9331,
    102.8667, 90.69854, 79.55382, 75.45756, 76.3409, 67.36531, 51.72295,
    50.51476, 47.67212, 46.14169, 43.00344, 41.73966, 40.72661, 38.58728,
    38.42667, 38.27389,
  97.91305, 89.27764, 77.35524, 71.30521, 73.60908, 74.77492, 77.46272,
    79.80039, 80.60065, 84.62599, 90.8973, 89.54195, 81.29315, 85.62866,
    87.70422, 89.70958, 95.6837, 99.76389, 95.67317, 83.48046, 64.30983,
    54.52576, 49.75257, 46.95249, 43.458, 41.5545, 40.4658, 38.96849,
    38.46059, 38.34632,
  90.6739, 83.49586, 71.47189, 66.29817, 69.63718, 72.00706, 73.61467,
    74.2882, 76.31255, 80.80669, 80, 68.95023, 68.2775, 67.59942, 67.45612,
    68.06652, 73.37462, 80.51225, 83.722, 82.01849, 74.06483, 63.52684,
    54.16888, 50.05524, 46.49297, 42.556, 40.72377, 39.17875, 38.44709,
    38.3654,
  86.08921, 78.91837, 69.57619, 65.33748, 66.91583, 67.3056, 67.03201,
    67.22113, 68.64203, 70.93098, 65.51932, 57.6067, 61.25626, 61.02438,
    59.412, 58.44392, 59.86541, 62.71836, 66.33434, 68.09883, 68.72127,
    68.82568, 62.64565, 55.42732, 49.28945, 43.96399, 40.76456, 39.2432,
    38.41924, 38.35968,
  89.91478, 82.71417, 73.93848, 69.33929, 69.28844, 64.92301, 64.37363,
    63.25104, 66.35577, 66.18214, 57.59477, 53.67617, 55.82885, 55.65163,
    54.8973, 54.72953, 54.28918, 55.22117, 57.94558, 59.60651, 60.56745,
    61.23742, 62.28148, 61.73995, 55.04165, 45.81582, 41.73833, 40.33367,
    38.72091, 38.31332,
  96.22019, 94.30519, 82.58127, 78.34268, 80.16803, 78.36786, 73.67401,
    68.86256, 68.24506, 64.87981, 58.16006, 58.6656, 59.7873, 60.26789,
    59.11499, 59.25807, 58.47302, 55.87978, 55.95253, 56.42534, 56.50771,
    56.57968, 56.28193, 58.40224, 59.4712, 52.02171, 44.8462, 42.94276,
    40.47649, 38.50661,
  103.1322, 101.9582, 94.86307, 92.4313, 91.52603, 88.29827, 89.72192,
    87.92863, 86.65819, 78.47902, 71.59839, 75.201, 75.50613, 76.8382,
    74.2476, 71.94089, 69.71259, 65.94781, 61.78626, 60.12468, 58.66825,
    57.49514, 56.53477, 56.26158, 58.3638, 58.98171, 53.04766, 45.68945,
    43.06419, 39.77514,
  101.5369, 99.32264, 85.49856, 83.27029, 83.84201, 83.05441, 82.92271,
    85.66534, 89.26856, 81.69162, 72.8013, 76.23702, 77.6788, 78.55439,
    77.41795, 76.41339, 73.09895, 70.28806, 67.00779, 63.5463, 61.45655,
    59.52782, 56.32794, 54.4483, 55.61762, 58.51554, 58.40624, 50.76715,
    45.69335, 42.11436,
  109.7399, 107.2637, 98.46599, 88.7953, 85.65356, 83.17748, 87.98727,
    91.85503, 87.02384, 79.82385, 79.55092, 80.78597, 81.83836, 80.27565,
    77.48136, 77.10548, 75.61158, 73.90582, 72.45335, 70.0526, 68.41711,
    66.30467, 61.8984, 58.58916, 58.81754, 59.70376, 60.16521, 53.00744,
    43.24108, 40.72552,
  112.7555, 109.3539, 97.95685, 89.13831, 84.27446, 80.83727, 85.92613,
    87.06067, 81.53278, 79.66013, 82.23614, 84.49486, 83.98357, 82.43639,
    80.10304, 78.10651, 76.20886, 75.1037, 74.41568, 73.32001, 73.22064,
    74.03725, 72.23831, 68.75835, 68.27646, 69.19231, 70.56777, 63.61987,
    47.08656, 39.00789,
  106.5682, 104.7169, 99.8156, 96.81371, 95.48809, 91.50829, 89.17104,
    83.93684, 76.91318, 78.62624, 79.47404, 79.60911, 81.02212, 79.62222,
    77.59593, 74.73975, 71.03423, 69.88772, 70.71247, 70.81953, 67.77856,
    63.62879, 59.89145, 59.20338, 60.93592, 62.86491, 64.20357, 66.19724,
    58.67926, 43.00834,
  83.46913, 84.68206, 88.89998, 92.63947, 96.74144, 99.02663, 91.11826,
    74.96637, 69.88091, 69.80641, 67.10819, 66.08418, 65.81705, 65.7931,
    65.39198, 63.52995, 61.00346, 59.61256, 56.89715, 53.72223, 52.6328,
    51.03465, 48.71298, 47.24392, 48.36881, 49.71294, 49.43232, 47.73986,
    48.21981, 44.3837,
  65.01742, 68.48584, 68.90866, 69.24368, 73.81794, 80.94191, 79.63815,
    66.01454, 59.20422, 62.65789, 64.2559, 65.93142, 65.62661, 62.73597,
    58.80689, 56.54796, 51.15404, 46.53704, 45.6589, 44.76653, 43.28651,
    43.59021, 43.66207, 43.64216, 44.02161, 45.012, 45.07114, 42.67548,
    40.19821, 38.30749,
  52.46587, 53.41888, 53.94504, 54.66728, 55.16697, 55.76105, 56.48406,
    57.20959, 57.97266, 58.96337, 60.5787, 60.68995, 57.90462, 57.48999,
    56.78829, 54.93846, 53.5454, 52.80107, 52.1042, 52.03443, 51.45575,
    49.35049, 49.21844, 50.89633, 51.85, 50.12283, 51.2252, 52.47503,
    42.34652, 38.63129,
  58.33091, 59.16814, 58.80792, 59.64523, 59.42625, 59.52033, 60.29508,
    61.08874, 62.006, 63.14038, 64.72884, 66.9458, 68.14115, 66.60711,
    65.48541, 65.17045, 63.61127, 63.7602, 64.09803, 64.51873, 64.1429,
    62.5945, 61.5325, 63.12758, 64.71585, 57.44534, 48.92653, 51.10071,
    42.86686, 39.60861,
  60.81027, 61.47013, 61.62665, 61.62085, 61.32498, 61.10899, 60.96418,
    61.04571, 61.17546, 61.23405, 61.61957, 62.7204, 63.87434, 65.2899,
    66.02633, 64.22383, 64.51958, 66.27862, 68.15726, 71.39606, 76.99988,
    81.83968, 81.87312, 79.09854, 74.987, 67.7557, 59.80035, 49.98306,
    42.31403, 40.12198,
  66.77396, 67.74462, 68.5826, 69.34888, 69.68853, 70.13744, 69.72043,
    68.8879, 68.72899, 68.26153, 67.32289, 66.98295, 65.82763, 64.17541,
    65.53214, 65.61134, 62.41877, 60.69698, 63.869, 67.97016, 74.13889,
    75.0746, 72.30746, 76.59286, 74.84041, 73.24091, 69.59689, 58.30151,
    46.3078, 39.61181,
  71.88238, 72.32327, 73.39684, 73.87787, 73.75562, 73.74304, 74.17983,
    73.93081, 74.86584, 75.49017, 75.59126, 77.95866, 78.95766, 77.34004,
    76.32442, 75.68729, 71.51793, 65.30631, 64.52087, 68.1445, 67.00458,
    59.10263, 60.79539, 66.56105, 71.35724, 72.21743, 72.01656, 77.89705,
    69.80515, 46.64268,
  76.65678, 79.575, 81.64473, 83.276, 81.92715, 81.54534, 84.02975, 83.75034,
    81.88835, 80.98206, 82.61867, 89.32891, 96.31886, 93.64616, 93.50824,
    94.55924, 91.49078, 83.27205, 73.04431, 69.81765, 62.53376, 54.94787,
    58.76851, 61.89058, 65.61664, 66.3795, 67.70316, 78.81903, 72.2793,
    43.03159,
  81.09195, 84.37225, 86.68777, 88.8675, 89.48571, 91.94321, 97.49734,
    101.4402, 99.50138, 93.90131, 88.11324, 78.19547, 67.97881, 67.91014,
    68.27054, 70.30219, 71.1105, 67.41386, 62.5611, 62.6415, 60.24426,
    59.09743, 61.12745, 64.44974, 64.56653, 61.22247, 64.93472, 71.10481,
    58.99749, 37.47754,
  82.05537, 84.46672, 86.93084, 89.22469, 90.40966, 95.86481, 98.15691,
    85.45131, 78.91667, 79.4789, 77.02123, 74.05607, 71.44606, 70.46711,
    69.13039, 68.86615, 70.03074, 68.45361, 63.96473, 62.67985, 62.87074,
    65.0433, 68.08757, 68.9679, 66.0871, 65.88314, 70.58997, 67.87531,
    51.78977, 38.16998,
  87.23768, 86.81514, 86.62732, 86.6622, 86.83162, 86.72679, 78.91789,
    79.00099, 81.48354, 82.53371, 83.39967, 83.46069, 83.85432, 88.55602,
    89.87321, 80.9726, 79.44797, 80.14142, 77.27541, 71.22643, 67.64635,
    71.40949, 76.35674, 74.60888, 69.54121, 74.31845, 73.19319, 59.50703,
    39.87627, 38.19049,
  110.2797, 108.9685, 100.4383, 97.63017, 96.44665, 87.47604, 72.36673,
    76.45721, 74.89281, 75.69225, 77.38181, 80.64272, 79.77558, 77.47653,
    75.67676, 79.49602, 80.46835, 79.55822, 77.44741, 76.65446, 77.46825,
    73.14168, 67.99011, 62.61248, 66.64644, 73.75414, 65.19688, 45.46327,
    37.87061, 36.73901,
  137.9318, 136.9127, 133.1569, 117.1013, 113.8155, 102.0478, 90.66288,
    88.99417, 88.60685, 83.83218, 73.18989, 61.72099, 59.3309, 59.23441,
    59.5097, 60.40184, 61.9553, 63.07303, 63.99577, 67.09175, 73.61337,
    70.33931, 60.28081, 59.05922, 63.00811, 60.26831, 46.73093, 38.55458,
    38.37391, 36.86341,
  145.4549, 142.8312, 144.5936, 143.4559, 139.8389, 113.47, 103.4282,
    93.22198, 86.0713, 80.00145, 74.61306, 70.54958, 71.62463, 70.22987,
    64.57471, 61.92139, 59.82952, 58.92164, 58.8398, 61.47328, 67.06215,
    65.15438, 58.19379, 64.98219, 67.4159, 53.84163, 39.92365, 42.52406,
    39.56823, 37.81379,
  141.1115, 142.952, 144.7579, 144.7977, 143.4815, 139.8222, 123.6979,
    109.8337, 112.1398, 101.025, 95.04625, 88.8387, 92.64529, 93.90467,
    82.66555, 68.18476, 67.79402, 65.88197, 63.78867, 64.65709, 64.75372,
    59.88062, 55.64145, 51.66223, 50.56941, 46.90009, 40.23331, 41.2091,
    40.75013, 38.6342,
  104.1494, 105.6943, 101.8838, 102.3385, 101.7232, 110.6317, 117.7878,
    117.2324, 104.7969, 106.746, 111.0634, 106.8255, 107.1721, 106.6829,
    98.33625, 81.98145, 73.66151, 76.66029, 77.76846, 71.02617, 61.81867,
    54.62453, 49.84725, 43.4001, 40.55854, 40.2954, 39.10053, 38.18819,
    38.57477, 38.03886,
  84.80904, 81.54189, 82.77512, 82.62403, 83.66985, 85.39481, 90.15256,
    88.60033, 84.73676, 84.48777, 80.89342, 77.49778, 80.33955, 84.80136,
    84.54022, 81.67938, 74.0424, 68.96289, 67.46188, 62.91584, 51.87022,
    50.04953, 44.55681, 42.40507, 41.77257, 40.73285, 39.45923, 38.33761,
    37.55909, 37.16238,
  87.00205, 89.20033, 89.33637, 88.56833, 86.98021, 88.1499, 89.8144,
    85.03209, 79.18732, 75.57057, 74.4741, 71.4671, 69.51859, 72.90327,
    69.86444, 68.20474, 67.31957, 60.98832, 57.54247, 52.98392, 46.23403,
    46.21449, 43.02368, 42.0535, 41.72431, 40.68594, 39.19373, 38.46092,
    37.76324, 37.19127,
  77.01357, 76.2759, 77.5259, 79.66513, 81.60023, 83.63052, 85.81748,
    87.68705, 85.97226, 82.45338, 78.40443, 83.04579, 87.39102, 81.72023,
    74.00305, 68.83765, 64.077, 60.17749, 58.0965, 53.59322, 45.82399,
    46.21906, 43.55527, 41.97024, 41.21893, 40.6129, 38.75433, 37.3703,
    37.2411, 37.07462,
  69.19201, 68.9774, 67.89189, 69.95579, 72.21719, 75.09203, 77.48955,
    79.70828, 81.55823, 82.02792, 87.78119, 92.35985, 90.36626, 89.28938,
    85.23027, 78.72182, 72.81857, 69.91591, 67.91461, 59.2271, 48.01296,
    45.77343, 43.86249, 42.61232, 40.5453, 39.67592, 38.72272, 37.10265,
    36.92637, 36.82603,
  74.65369, 68.07811, 60.23028, 56.97057, 59.38233, 60.3961, 62.28905,
    64.05864, 64.41704, 66.86732, 70.52318, 69.39232, 65.40941, 67.81727,
    69.21756, 72.17949, 77.88602, 82.0509, 79.94831, 71.10511, 57.86733,
    49.61034, 45.70458, 43.80373, 41.18448, 39.6352, 38.6389, 37.36745,
    36.95043, 36.86007,
  70.51161, 65.62608, 57.60493, 53.33158, 55.01476, 55.98705, 57.39352,
    58.94621, 61.18125, 65.09421, 64.61839, 58.26908, 57.93584, 56.64238,
    55.72073, 56.21814, 59.84291, 65.03311, 67.46912, 67.08951, 62.50233,
    55.69767, 49.01612, 45.84238, 43.21478, 40.39547, 38.86257, 37.53509,
    36.93986, 36.86757,
  73.00435, 68.38608, 59.78244, 55.4476, 55.77061, 55.90837, 56.74266,
    58.04147, 60.22324, 62.03082, 58.70448, 54.88682, 57.20851, 56.13334,
    54.42349, 53.51408, 54.03176, 55.33623, 56.94226, 57.14455, 57.81321,
    58.09971, 53.95632, 49.64056, 45.28997, 41.44526, 38.91734, 37.61313,
    36.96705, 36.88477,
  81.09018, 77.58298, 68.98744, 65.41644, 64.92265, 62.45295, 61.99505,
    61.66154, 63.50715, 63.20453, 58.04159, 55.20718, 56.18386, 55.56283,
    54.19532, 53.60757, 52.48278, 52.141, 53.13055, 53.42852, 53.09167,
    52.99956, 53.71776, 53.06214, 49.10925, 42.83966, 39.71127, 38.45586,
    37.25366, 36.89216,
  88.39966, 88.67001, 79.50238, 76.46262, 78.06461, 77.13921, 74.47072,
    70.75746, 70.25475, 67.6254, 62.48842, 62.53325, 62.18389, 61.2349,
    59.21134, 58.352, 56.68169, 53.77056, 52.61003, 51.96907, 51.03787,
    50.0964, 49.43531, 50.97231, 51.95366, 46.99427, 41.90151, 40.30129,
    38.51826, 37.0482,
  91.18521, 90.84029, 85.33226, 83.69388, 83.86301, 82.23652, 81.9923,
    80.88201, 82.19736, 77.00401, 71.40675, 72.68298, 73.21935, 72.91242,
    69.97812, 67.26003, 64.48759, 60.64653, 57.00735, 54.97987, 52.78127,
    50.89349, 49.78268, 49.48815, 51.03023, 51.36597, 47.20507, 42.06394,
    40.11972, 37.91311,
  92.6696, 88.75754, 80.71476, 77.81867, 77.66256, 76.4693, 77.34325,
    80.87939, 84.79137, 79.23787, 72.67897, 73.66005, 74.11346, 74.03613,
    72.22073, 70.14471, 66.56641, 63.39877, 60.4497, 57.56728, 55.39392,
    52.86035, 50.03714, 48.4991, 49.36648, 51.20061, 50.68643, 45.07333,
    41.652, 39.30273,
  94.41593, 91.81048, 84.57076, 78.4229, 75.14491, 73.59993, 77.18072,
    81.42626, 80.30359, 74.76689, 73.81738, 74.24688, 74.57352, 72.94358,
    70.4901, 69.1636, 67.04447, 64.79598, 63.16405, 61.08677, 59.96649,
    58.36488, 54.72206, 51.91859, 51.91138, 52.25107, 52.16977, 46.67983,
    40.19328, 38.42542,
  90.26989, 86.84029, 79.2751, 74.30704, 70.49265, 66.90875, 70.00555,
    70.97631, 68.72115, 66.66523, 68.03282, 68.99155, 69.53672, 68.73626,
    67.38521, 65.83488, 63.98537, 62.63925, 61.91385, 60.73946, 60.5345,
    61.24974, 59.94096, 57.50032, 57.33199, 58.12906, 58.95367, 53.6182,
    42.58307, 37.39094,
  79.2665, 77.61841, 74.91779, 73.51118, 72.58127, 68.24789, 65.71275,
    62.35065, 57.92133, 58.66721, 59.27168, 60.4325, 61.65257, 62.31686,
    62.02885, 60.89756, 59.04785, 57.94907, 58.37868, 58.29873, 56.45464,
    53.90053, 51.42536, 50.62939, 51.6433, 52.80801, 53.54841, 54.60319,
    49.87688, 39.95182,
  60.53939, 60.53329, 62.21102, 64.22414, 66.79552, 68.54858, 63.39817,
    54.58982, 51.60409, 52.50725, 52.00461, 52.0815, 52.61569, 52.80509,
    52.58696, 52.51948, 51.35854, 50.39452, 48.90084, 47.26087, 46.52775,
    45.77876, 44.4952, 43.45982, 44.08308, 44.72377, 44.12904, 42.83836,
    43.42281, 40.82054,
  49.86558, 50.4029, 50.23647, 49.69782, 52.10847, 56.8567, 57.36614,
    49.22219, 45.812, 48.14127, 49.85447, 51.32222, 51.32268, 49.69947,
    47.78737, 47.00845, 44.25819, 41.5532, 41.23651, 40.73722, 39.87369,
    40.28107, 40.67064, 40.87915, 41.00065, 41.44424, 41.20728, 39.71503,
    38.27743, 36.9224,
  47.52715, 47.71143, 47.69094, 47.70519, 47.60329, 47.65314, 47.72752,
    47.81694, 47.99063, 48.33658, 49.14524, 48.99542, 46.95399, 47.01431,
    46.73027, 45.60438, 45.0751, 45.05522, 45.06873, 45.61126, 45.67648,
    44.40953, 44.88531, 46.82147, 48.05681, 47.1992, 48.50003, 49.55259,
    40.34058, 37.01073,
  53.39607, 53.75097, 53.12675, 53.58266, 53.23701, 53.14809, 53.58467,
    54.00821, 54.61561, 55.29443, 56.1907, 57.38311, 57.86861, 56.36432,
    55.13549, 54.83661, 53.64799, 53.9064, 54.47691, 54.90578, 54.50041,
    53.67144, 53.81453, 56.43047, 58.7233, 53.12935, 45.22474, 48.19734,
    40.52012, 37.75874,
  54.25436, 54.36491, 54.18785, 54.11533, 53.99686, 54.0744, 54.35406,
    54.85448, 55.63716, 56.44633, 57.33511, 58.63823, 59.91836, 61.18517,
    61.6361, 59.98911, 60.36887, 61.91264, 63.62688, 66.38683, 71.3226,
    75.79812, 75.22135, 71.05033, 66.67975, 61.19157, 54.5397, 46.85723,
    40.2562, 38.40195,
  58.61281, 58.76453, 58.97925, 59.2758, 59.24321, 59.42374, 59.20222,
    58.68357, 58.85999, 59.07659, 58.91913, 59.47304, 59.61474, 59.29127,
    61.28605, 62.04733, 60.03065, 59.25425, 62.33583, 65.97884, 71.8584,
    72.28049, 66.60088, 69.10594, 66.36426, 64.37833, 62.64557, 52.25597,
    42.32909, 37.63998,
  64.09219, 63.92905, 64.5066, 64.73837, 64.45662, 64.09351, 64.26305,
    64.21625, 65.12435, 65.4867, 65.10611, 66.60521, 67.41293, 66.91056,
    67.20838, 67.15768, 64.62285, 61.40824, 62.2817, 66.22995, 66.02799,
    57.95618, 58.70641, 62.74063, 66.05869, 66.80038, 64.70963, 69.36674,
    64.10676, 45.06465,
  68.53807, 70.45395, 72.00331, 73.37212, 72.34535, 72.05636, 74.43736,
    74.85048, 74.53233, 75.30042, 77.71658, 84.07738, 90.03934, 87.34523,
    87.19262, 87.14584, 85.71584, 78.74896, 69.58612, 66.55556, 59.2418,
    52.46512, 56.36904, 59.1412, 62.33493, 62.96472, 63.42983, 72.78054,
    67.9731, 41.70397,
  70.67447, 73.01537, 74.76366, 76.47151, 76.87609, 79.21681, 85.21472,
    89.90936, 88.85316, 84.28622, 79.55106, 70.75363, 61.56597, 62.08443,
    62.73693, 64.13754, 64.52668, 61.80832, 57.79391, 57.3896, 54.9376,
    53.71417, 56.10531, 59.34422, 59.9981, 57.76738, 60.818, 66.47707,
    57.07457, 35.96701,
  70.71736, 73.2198, 75.4544, 77.64544, 78.76483, 83.51671, 85.77644,
    73.20757, 66.2672, 66.6089, 64.31536, 61.74875, 59.91144, 59.82748,
    59.61313, 60.40895, 62.06231, 61.04195, 57.73304, 57.22284, 57.27258,
    58.83143, 61.53003, 62.81305, 60.6636, 61.32609, 67.0481, 65.02597,
    49.25213, 36.39582,
  75.04578, 76.05849, 76.85171, 77.83107, 78.81485, 79.55145, 71.95092,
    71.34247, 73.27493, 73.59225, 73.99069, 73.78468, 74.18898, 78.34731,
    79.53413, 72.15236, 71.01752, 71.54427, 69.77425, 65.14603, 62.54216,
    65.94527, 70.11693, 68.74657, 63.87117, 68.13873, 68.89942, 57.579,
    38.13071, 36.67639,
  90.82432, 91.22819, 84.11928, 83.01658, 83.65078, 77.32457, 64.07585,
    69.02879, 68.32568, 69.57291, 71.53667, 74.87287, 73.78365, 72.33682,
    70.4178, 73.19534, 73.92063, 72.69841, 70.57416, 69.62349, 70.39189,
    67.32897, 63.24133, 58.7964, 62.65533, 70.13368, 62.97272, 43.91114,
    36.20945, 35.40004,
  121.7358, 115.5963, 108.941, 94.8515, 94.32858, 84.48852, 75.06284,
    75.39836, 75.92599, 72.86716, 65.07489, 55.64188, 54.78237, 54.94764,
    55.13922, 56.41941, 57.98217, 58.6914, 59.1001, 61.43049, 66.94228,
    64.68069, 56.15011, 54.91618, 58.98324, 57.26005, 44.86809, 36.35097,
    36.75741, 35.46938,
  130.0083, 125.9778, 126.4418, 125.5933, 117.8493, 93.83056, 85.72549,
    76.88536, 70.53762, 66.92058, 63.21043, 60.82874, 61.82048, 60.83408,
    57.35813, 55.77104, 54.86322, 54.58794, 54.93271, 57.32164, 62.59848,
    61.92276, 56.08369, 62.096, 64.43832, 51.80509, 37.41121, 40.04517,
    37.54396, 36.252,
  129.3634, 129.6852, 130.5781, 130.1695, 128.5608, 124.4086, 106.9369,
    89.42825, 95.27291, 84.94197, 80.86372, 76.57815, 80.10724, 81.50221,
    72.14244, 59.63489, 60.13273, 59.18481, 58.12424, 59.36161, 60.5181,
    57.50486, 53.97092, 50.69368, 49.58999, 45.20227, 38.54151, 39.51013,
    38.85051, 37.0805,
  100.4761, 101.8055, 97.76882, 97.51513, 94.97039, 100.1563, 105.1073,
    105.4721, 93.90475, 95.05702, 100.2522, 96.32455, 95.87425, 95.44616,
    87.6059, 72.89488, 66.71802, 69.80849, 71.35411, 65.37546, 57.16652,
    50.98716, 47.15959, 41.39916, 38.61449, 38.5075, 37.34921, 36.67897,
    36.91942, 36.51962,
  75.39845, 72.00202, 73.56777, 73.67051, 74.58586, 75.87909, 79.57819,
    79.59557, 76.38321, 77.01397, 74.3998, 71.54858, 73.78055, 77.15332,
    76.27089, 75.15325, 67.44357, 63.34839, 61.97748, 58.3194, 48.45586,
    46.69215, 41.53877, 39.70643, 39.40318, 38.55982, 37.48477, 36.57436,
    36.00772, 35.7276,
  74.22621, 76.1967, 76.18312, 75.0762, 73.07559, 73.80676, 75.10828,
    71.43681, 67.03303, 64.34844, 64.31221, 61.90576, 60.895, 64.52055,
    62.42281, 60.74152, 60.78197, 55.75508, 53.15733, 49.46642, 43.13844,
    43.26804, 40.5036, 39.5852, 39.37218, 38.63546, 37.46, 36.80083,
    36.20235, 35.76896,
  67.2812, 66.76433, 67.40529, 68.65012, 69.49551, 69.9513, 70.94183,
    72.55388, 71.10865, 68.11987, 64.48709, 68.09137, 71.90413, 67.9155,
    62.58765, 59.16528, 56.00327, 53.11778, 52.19121, 49.51062, 43.17977,
    43.63518, 41.19363, 39.64804, 39.00138, 38.60329, 37.13008, 36.00742,
    35.78788, 35.64145,
  62.01679, 62.55573, 61.83398, 63.51104, 65.24012, 66.95038, 68.43759,
    70.33508, 71.8735, 71.71974, 75.42384, 78.50363, 77.13043, 76.02556,
    71.39039, 66.4583, 61.41263, 59.17544, 58.29893, 52.99265, 44.47844,
    42.9276, 41.15416, 40.08474, 38.48576, 37.81678, 37.09546, 35.72623,
    35.51723, 35.44556,
  69.01489, 63.9236, 56.91918, 54.02032, 56.28794, 57.18936, 58.70985,
    60.25361, 60.76468, 62.74603, 66.00085, 65.28656, 61.29754, 62.75529,
    63.62498, 65.72498, 70.08767, 73.18571, 70.95476, 63.91636, 52.68092,
    45.79595, 42.34283, 40.92082, 39.10669, 37.90332, 37.04688, 35.91135,
    35.52809, 35.47698,
  66.29507, 61.4434, 54.30882, 50.12144, 51.49212, 52.10635, 53.06798,
    54.07692, 55.74458, 58.98917, 59.1507, 54.21179, 54.10165, 53.15389,
    52.45797, 52.76702, 55.65142, 59.84153, 61.69853, 60.82777, 56.23957,
    50.40459, 44.9134, 42.46748, 40.68672, 38.51518, 37.29436, 36.11228,
    35.51453, 35.48865,
  66.41719, 61.77589, 53.81147, 49.52716, 49.73048, 49.83093, 50.31675,
    51.06039, 52.69405, 54.41653, 52.3323, 49.31866, 51.37787, 50.7449,
    49.408, 48.70271, 49.31282, 50.66795, 52.11094, 51.87625, 51.56592,
    51.51987, 48.681, 45.23353, 42.08648, 39.25251, 37.33391, 36.16447,
    35.57184, 35.50702,
  70.75359, 67.00508, 58.85008, 54.79897, 54.3317, 52.39641, 52.16833,
    51.93204, 53.48775, 53.68922, 49.90919, 47.87569, 48.98927, 48.74102,
    47.99459, 47.86335, 47.40487, 47.51397, 48.26948, 48.23637, 48.02231,
    48.09286, 48.41598, 47.82694, 44.42292, 40.04814, 37.79257, 36.70959,
    35.77388, 35.51952,
  76.73022, 75.58748, 66.98538, 63.40252, 64.2645, 63.26393, 61.26039,
    58.50153, 58.24721, 56.42084, 52.27414, 52.34974, 52.42907, 52.06213,
    50.87347, 50.60867, 49.84934, 47.98499, 47.33717, 46.93518, 46.36227,
    45.97939, 45.46433, 46.15676, 46.4583, 42.76997, 39.29367, 38.10838,
    36.74297, 35.62788,
  79.84322, 79.08946, 73.49928, 71.21352, 70.76851, 69.22945, 69.15942,
    68.27425, 69.54953, 65.8889, 61.32281, 62.55004, 63.37095, 63.1978,
    61.05264, 58.98702, 56.97582, 54.29316, 51.59217, 50.06768, 48.62111,
    47.31696, 46.29536, 45.59639, 46.46212, 46.70548, 43.6252, 39.46025,
    37.99401, 36.28297,
  79.62987, 75.19214, 69.03517, 66.43625, 66.47305, 65.67154, 66.46368,
    69.43311, 72.87868, 68.63898, 63.28314, 64.23787, 64.85999, 65.28198,
    64.09408, 62.81519, 60.31917, 57.69461, 54.85205, 52.49395, 51.12257,
    49.21563, 46.74266, 45.2207, 45.87414, 47.37465, 46.95618, 42.42127,
    39.5306, 37.51346,
  80.86629, 77.76277, 72.45614, 67.8425, 65.96096, 65.23403, 68.19216,
    71.86085, 71.48067, 66.98257, 66.00571, 66.29941, 66.76088, 66.17136,
    64.33129, 63.16341, 61.68631, 59.8221, 57.57319, 55.58382, 54.90349,
    53.32061, 49.61161, 46.95433, 46.99669, 47.5629, 47.82611, 43.61737,
    38.3674, 36.78845,
  78.86295, 75.07961, 69.83606, 66.01949, 63.99257, 62.22763, 65.15112,
    66.2855, 64.83798, 63.21317, 64.29394, 64.90594, 65.51062, 65.2748,
    64.14604, 62.67532, 61.73047, 60.9098, 59.32258, 57.98319, 58.3912,
    58.79079, 56.53105, 53.54525, 52.64767, 53.33434, 53.96669, 49.31364,
    39.86719, 35.85355,
  72.15046, 70.79408, 67.35577, 65.82154, 65.78777, 63.66013, 62.21133,
    59.80919, 56.84158, 57.40907, 58.04926, 58.99635, 60.2893, 61.10316,
    60.68317, 59.3865, 58.04659, 57.64049, 57.17659, 56.66227, 55.55767,
    53.65234, 51.25917, 50.01657, 50.33763, 50.90582, 51.13012, 51.17599,
    46.37868, 37.85629,
  57.95638, 58.61849, 59.34864, 60.10465, 61.90224, 63.60062, 59.83956,
    52.76663, 50.5782, 51.16177, 50.56899, 50.52261, 51.11183, 51.53503,
    51.61509, 51.39952, 50.50672, 49.84277, 48.22515, 46.39981, 45.46767,
    44.66545, 43.70125, 42.97421, 43.32386, 43.61817, 42.8899, 41.39594,
    41.23526, 38.90569,
  48.8336, 49.58933, 49.65432, 49.21402, 51.00608, 54.8737, 55.21846,
    48.61511, 45.82269, 47.73381, 48.88345, 49.92965, 49.84351, 48.30417,
    46.5766, 45.6039, 43.04562, 40.98045, 40.68615, 40.03383, 39.10166,
    39.4108, 39.88882, 40.05337, 40.0172, 40.19024, 39.76172, 38.28977,
    36.87894, 35.58818,
  38.3594, 38.48664, 38.68625, 38.85381, 38.93841, 39.04752, 39.15026,
    39.3515, 39.74475, 40.32053, 41.30537, 41.34294, 39.75102, 40.20748,
    40.38564, 40.00824, 40.12056, 40.59447, 41.21729, 42.19416, 42.65512,
    42.0204, 42.57635, 44.16167, 45.61368, 45.87206, 47.42202, 48.47037,
    41.47346, 38.96743,
  41.27598, 41.50602, 41.33658, 41.80527, 41.54796, 41.39154, 41.59109,
    41.84231, 42.21607, 42.70283, 43.3847, 44.25095, 44.66998, 43.68916,
    43.17867, 43.69318, 43.32583, 44.24296, 45.525, 46.66071, 47.07705,
    47.42816, 49.05431, 52.78249, 56.00026, 51.89018, 45.34689, 48.14504,
    41.98094, 39.59628,
  44.33008, 44.48875, 44.62408, 44.75868, 44.78112, 44.90639, 45.11568,
    45.49269, 46.00784, 46.54791, 47.29322, 48.46709, 49.5604, 50.72178,
    51.53188, 51.04919, 52.32711, 54.47438, 56.7413, 60.09805, 65.23173,
    70.65634, 71.43712, 67.88353, 64.10852, 58.88958, 53.6677, 47.53813,
    41.89719, 40.27485,
  48.65215, 49.39333, 50.19327, 51.03858, 51.54211, 52.09579, 52.16092,
    52.1258, 52.61034, 53.28671, 53.71058, 54.60896, 55.25143, 55.46864,
    57.60534, 59.06254, 58.52416, 58.71382, 62.2531, 66.48186, 72.13275,
    71.76151, 65.28241, 66.29902, 62.54203, 61.02502, 59.418, 50.69614,
    42.29019, 39.25853,
  51.41176, 51.25776, 51.96007, 52.38184, 52.41179, 52.26483, 52.50635,
    52.73804, 53.63855, 54.23775, 54.1853, 55.34588, 56.61173, 57.65345,
    59.0335, 60.71741, 60.57743, 59.82684, 62.61525, 67.25323, 66.69028,
    58.57806, 57.68939, 61.4199, 63.76377, 63.73757, 62.55925, 67.54815,
    63.10444, 46.48344,
  54.79307, 56.35385, 58.102, 59.85814, 59.83598, 60.61227, 63.67981,
    65.50556, 67.33312, 70.42491, 75.31592, 84.18758, 91.9418, 89.36871,
    89.71198, 90.88312, 88.07919, 81.38634, 73.89299, 70.43857, 62.76228,
    55.23664, 59.43716, 62.21561, 65.37212, 66.02925, 67.21336, 76.77554,
    70.96632, 43.81834,
  64.0258, 67.57359, 70.71793, 74.04998, 76.39859, 80.97263, 89.57381,
    96.58604, 96.09054, 91.6553, 88.30258, 80.49078, 70.93723, 70.42391,
    70.41943, 70.91695, 69.92493, 65.66424, 60.96693, 59.85569, 56.75843,
    55.31541, 57.91361, 60.99332, 61.71172, 60.10799, 63.86219, 69.6624,
    58.8764, 38.11148,
  67.5802, 70.60153, 73.21455, 75.93548, 77.53546, 82.69812, 84.82276,
    70.56587, 62.19547, 61.51499, 58.19049, 54.8675, 52.73676, 53.03553,
    53.84785, 55.65405, 56.97686, 56.32427, 54.42665, 54.72652, 54.97677,
    56.34488, 59.17311, 61.21238, 60.29735, 61.6419, 67.50206, 66.0562,
    51.61517, 38.18664,
  68.16219, 69.35635, 70.2468, 70.85155, 72.13375, 72.05611, 62.45279,
    59.67043, 60.93887, 60.94373, 61.27613, 61.56585, 62.97341, 67.10892,
    68.99905, 63.89137, 64.34984, 66.08266, 65.63176, 62.74624, 61.2968,
    65.09399, 69.03314, 68.02651, 64.3107, 68.9444, 69.98431, 59.14256,
    40.25044, 38.8345,
  75.20155, 78.53009, 75.55286, 76.77025, 78.50563, 73.16853, 60.38304,
    66.0621, 66.74426, 69.38081, 71.91315, 75.43316, 75.57583, 74.28115,
    72.30139, 74.17251, 74.89745, 73.991, 72.33401, 71.90291, 72.64556,
    70.28772, 66.89291, 62.71478, 66.12096, 72.74539, 66.04765, 46.14257,
    38.19526, 37.82,
  79.06432, 79.22083, 80.51353, 80.03922, 83.01392, 77.5993, 70.47061,
    73.69833, 75.77318, 73.90322, 66.96317, 58.91482, 58.08069, 58.86291,
    59.06271, 59.97591, 61.2627, 61.72344, 62.06807, 64.42113, 69.11852,
    66.55734, 58.6877, 57.80341, 62.64282, 61.12867, 47.64565, 38.26732,
    38.83613, 37.78957,
  99.31726, 91.82668, 97.24818, 98.09219, 90.44119, 76.52396, 76.06886,
    68.58612, 62.82335, 61.36733, 57.80708, 56.36752, 58.20745, 58.00779,
    56.31874, 56.10012, 55.44136, 55.851, 56.49156, 58.97575, 64.07895,
    63.84384, 59.27187, 65.11703, 66.46178, 53.46832, 38.97547, 41.29328,
    39.27301, 38.34888,
  118.7949, 120.2063, 121.2741, 120.1825, 117.3903, 112.5634, 89.65865,
    75.47024, 81.88712, 72.51256, 68.70677, 66.2389, 70.11572, 71.85285,
    66.05868, 56.63152, 57.79242, 57.86455, 58.22467, 60.43764, 63.11293,
    62.15231, 59.46388, 55.84974, 53.3857, 47.45913, 40.30969, 41.5089,
    40.5299, 39.14387,
  113.1194, 112.8151, 111.6953, 109.0224, 104.6301, 104.7408, 105.3922,
    104.6216, 91.59235, 91.4066, 95.30145, 91.88469, 89.35066, 88.65408,
    82.21065, 69.88592, 66.44732, 70.57354, 72.5535, 66.82298, 60.29974,
    55.22295, 50.49913, 44.74664, 41.48107, 40.99723, 39.84999, 39.24151,
    39.28164, 38.8133,
  87.25065, 82.08812, 82.60198, 81.62447, 81.98558, 84.18254, 87.73021,
    85.12424, 80.66867, 80.00032, 77.40102, 74.66609, 75.86411, 77.939,
    77.0674, 76.12827, 70.04117, 65.84746, 64.29522, 59.9884, 50.89949,
    48.49249, 43.54397, 41.17884, 41.0837, 40.52081, 39.63127, 38.8086,
    38.36597, 38.09693,
  72.54544, 73.77015, 73.97282, 73.02431, 71.55222, 71.90727, 72.99271,
    70.33289, 66.19935, 63.96632, 63.64045, 61.72627, 61.35807, 64.27918,
    62.24828, 61.28819, 61.10764, 56.25852, 53.94131, 50.10638, 44.51864,
    44.52237, 41.81869, 41.07228, 41.04861, 40.57637, 39.67775, 39.06948,
    38.46741, 38.06771,
  61.72338, 60.30972, 60.41996, 61.0494, 61.66001, 61.97306, 62.37948,
    63.30938, 62.60282, 60.75793, 58.05845, 61.11972, 65.09897, 62.55997,
    58.66087, 56.42375, 54.40133, 52.55084, 52.21503, 49.98676, 44.56701,
    44.79099, 42.42629, 41.19668, 40.90337, 40.65873, 39.38583, 38.39596,
    38.11766, 37.9896,
  57.82093, 58.30208, 57.56561, 58.39499, 59.0837, 59.91694, 60.66845,
    61.92613, 62.94035, 62.36153, 65.13193, 67.6041, 66.47717, 65.52087,
    61.94701, 57.61194, 54.0597, 53.48663, 54.48555, 51.22029, 44.82753,
    43.95235, 42.39185, 41.55842, 40.40103, 39.96492, 39.25957, 38.09782,
    37.85984, 37.79822,
  68.64328, 63.92284, 57.24426, 53.8134, 55.1246, 55.13439, 55.91553,
    56.91897, 56.97878, 58.43526, 61.1162, 60.50806, 57.13112, 58.1827,
    58.24335, 59.96355, 64.49158, 68.157, 66.90421, 60.97125, 51.76606,
    46.30312, 43.57954, 42.52242, 41.02728, 40.11295, 39.29933, 38.23853,
    37.84486, 37.80551,
  66.30045, 61.92465, 55.22651, 51.4432, 52.74202, 53.17375, 54.05547,
    55.14965, 56.82805, 59.71462, 60.17316, 56.3906, 56.45501, 55.77498,
    55.02813, 55.461, 58.12075, 61.56245, 62.26125, 60.30584, 55.13134,
    49.74449, 45.58523, 43.99998, 42.43298, 40.61242, 39.52522, 38.37178,
    37.82684, 37.82893,
  63.18811, 59.40529, 52.70387, 49.46875, 50.4016, 50.87206, 51.60379,
    52.53667, 54.1479, 55.79179, 54.13697, 51.59267, 53.37613, 52.77108,
    51.43233, 50.8016, 51.40388, 52.4806, 53.28821, 52.49354, 51.7295,
    51.11102, 48.49039, 46.079, 43.68397, 41.31731, 39.47316, 38.40894,
    37.88879, 37.85415,
  61.86515, 58.81199, 52.05971, 48.96988, 49.44485, 48.66768, 49.26654,
    49.70033, 51.43773, 51.72206, 48.64756, 47.26199, 48.52612, 48.51771,
    47.98618, 48.07103, 48.10479, 48.54401, 49.29953, 49.38497, 49.14136,
    48.73056, 48.65409, 47.91444, 45.40678, 41.75961, 39.72815, 38.71912,
    38.01918, 37.87624,
  62.7821, 61.44529, 53.9785, 51.06473, 52.58657, 52.32045, 51.35744,
    49.72314, 49.86963, 48.84758, 46.11668, 46.72654, 47.52589, 48.00689,
    47.85763, 48.33217, 48.40733, 47.46996, 47.3786, 47.34686, 47.01484,
    46.51315, 45.95634, 46.59649, 46.86558, 43.57175, 40.71659, 39.83173,
    38.73212, 37.94619,
  68.74124, 68.05402, 62.89931, 60.8579, 60.69193, 59.18029, 59.20206,
    58.79541, 60.32124, 58.09826, 55.22609, 57.05676, 58.29109, 58.77959,
    57.54306, 56.40703, 55.29413, 53.27814, 51.2733, 50.0891, 48.84554,
    47.92871, 47.04419, 46.55239, 47.30445, 47.14655, 44.31329, 40.92695,
    39.72704, 38.44151,
  70.89504, 67.19599, 61.51067, 59.24704, 59.25144, 58.41502, 59.29379,
    62.25089, 65.86737, 63.0744, 59.15462, 60.66122, 61.86865, 62.71132,
    61.70822, 60.82412, 59.16349, 57.36784, 55.2059, 53.22257, 51.83596,
    50.23922, 47.99324, 46.62446, 47.26675, 48.23378, 47.57511, 43.64622,
    41.20182, 39.61893,
  73.46346, 70.83692, 65.83082, 61.79086, 60.48131, 59.87132, 62.65198,
    66.31635, 66.55135, 62.92915, 62.15436, 62.80284, 63.74432, 63.45297,
    61.57546, 60.85023, 59.82583, 58.28684, 56.53584, 54.91762, 53.90218,
    52.33736, 49.14314, 47.20258, 47.24704, 47.32636, 47.5672, 44.64436,
    40.47714, 39.18925,
  74.77485, 71.41239, 66.49354, 62.80729, 61.48551, 60.18919, 63.11134,
    64.88857, 63.94073, 62.33352, 63.28998, 63.82739, 64.30762, 64.00505,
    62.71139, 62.02155, 61.39256, 60.39151, 58.82524, 57.69627, 57.77391,
    57.62581, 55.68266, 53.06247, 51.77673, 51.07251, 51.08871, 48.01861,
    41.26834, 38.31995,
  73.44793, 71.14986, 67.8118, 66.7153, 67.078, 65.71835, 65.15335, 63.81404,
    61.59122, 62.06841, 62.8283, 63.56386, 64.6795, 65.21382, 64.40112,
    63.36454, 62.17961, 61.26448, 60.46854, 59.98513, 58.6085, 56.24437,
    53.53759, 52.15398, 51.80547, 51.18317, 50.47272, 50.10918, 46.38468,
    39.77057,
  60.44284, 60.68675, 61.54242, 62.18796, 63.90266, 65.22615, 62.16258,
    56.47998, 54.74208, 55.12955, 54.84048, 54.98063, 55.69656, 56.45095,
    56.64172, 56.57781, 55.84702, 54.6885, 52.62006, 50.89586, 49.93447,
    48.61407, 47.11548, 46.20334, 46.21129, 45.90716, 44.88933, 43.50583,
    43.02877, 40.78374,
  54.98767, 55.4254, 55.85916, 55.59505, 57.4294, 60.93606, 60.93008,
    54.7672, 52.25771, 53.94656, 55.01315, 55.65344, 55.16274, 53.44658,
    51.60811, 50.46987, 47.98755, 45.82291, 45.18692, 44.33467, 43.41838,
    43.4888, 43.63709, 43.60773, 43.37589, 43.05869, 42.15627, 40.61737,
    39.26148, 38.03553,
  33.98166, 34.00969, 34.10328, 34.15559, 34.20912, 34.29912, 34.33254,
    34.402, 34.55615, 34.92081, 35.64183, 35.64775, 34.60037, 34.91926,
    35.01191, 34.65622, 34.58357, 34.7167, 34.96252, 35.54719, 35.76565,
    35.30959, 35.65049, 36.8679, 38.38026, 39.02265, 40.37909, 41.18304,
    36.378, 34.67983,
  34.88897, 35.0327, 34.91041, 35.26147, 35.1781, 35.15928, 35.29407,
    35.46518, 35.72619, 36.05968, 36.50871, 37.02468, 37.22649, 36.47961,
    35.93125, 36.00354, 35.40109, 35.76191, 36.41056, 37.08376, 37.38171,
    38.02262, 40.17242, 44.47586, 48.34136, 44.98656, 39.39031, 41.57857,
    36.98275, 35.15961,
  35.34279, 35.30275, 35.34188, 35.41005, 35.42601, 35.57901, 35.76849,
    36.01913, 36.31742, 36.63676, 37.06945, 37.75757, 38.38617, 39.00566,
    39.29712, 38.89432, 39.81488, 41.5451, 43.6262, 47.0329, 52.51432,
    58.95256, 61.23259, 59.09075, 56.25217, 51.42072, 46.96254, 41.1864,
    36.93851, 35.73152,
  36.34928, 36.71658, 37.41472, 38.30659, 39.19822, 40.15119, 40.58348,
    40.84547, 41.41839, 42.02724, 42.43242, 43.28026, 43.954, 44.22783,
    46.25352, 48.21084, 48.81926, 50.19585, 54.28822, 59.39486, 65.63922,
    65.32294, 58.87175, 58.0959, 53.80462, 53.19566, 52.04446, 43.96078,
    36.59348, 34.82388,
  39.95188, 40.5337, 41.72209, 42.81274, 43.47403, 43.73966, 43.78314,
    43.43525, 43.43072, 43.25241, 43.0405, 44.17677, 45.93773, 47.95831,
    50.34047, 53.06017, 54.21248, 54.65882, 57.90076, 62.1534, 60.78767,
    52.16764, 49.75038, 52.58489, 54.20932, 54.72909, 54.97567, 60.24065,
    56.71322, 41.79917,
  42.4273, 43.19513, 43.98682, 44.55588, 43.8477, 43.53033, 44.89177,
    46.24355, 48.70422, 52.87334, 59.30121, 70.36674, 80.09968, 79.18651,
    80.38411, 81.64536, 79.25523, 74.41807, 67.79875, 63.52172, 55.32954,
    47.60529, 51.82439, 54.55497, 57.83564, 59.45903, 61.64112, 71.8107,
    66.57297, 40.17957,
  44.51137, 46.22844, 48.44579, 51.30885, 54.42662, 60.70291, 72.07384,
    83.27184, 87.50628, 87.78787, 88.95121, 84.99555, 77.11046, 76.00713,
    74.82414, 73.49837, 71.18484, 64.8028, 58.13859, 55.82105, 52.02531,
    50.69549, 53.68095, 56.38686, 57.34072, 56.71807, 60.98373, 66.66195,
    54.55928, 34.06287,
  53.69935, 58.90457, 64.33008, 70.72495, 76.88264, 87.1782, 93.971,
    83.37119, 75.95799, 74.00674, 69.16064, 63.43948, 58.94361, 57.26529,
    55.97991, 55.83708, 55.2733, 53.01321, 50.44027, 50.20121, 49.98844,
    50.84635, 53.23079, 55.1944, 54.91931, 56.67214, 62.91391, 61.98973,
    46.90763, 34.01427,
  66.49007, 71.38322, 74.79462, 77.66198, 80.67655, 80.47552, 69.39317,
    62.77628, 61.1567, 58.62948, 56.47977, 55.23641, 55.68604, 58.47354,
    59.42731, 55.39167, 55.56084, 56.82399, 56.22384, 54.03913, 52.90763,
    55.91472, 59.88388, 59.93683, 58.26493, 64.11914, 67.44514, 56.36761,
    36.02909, 34.54762,
  73.19537, 76.24374, 73.76402, 73.94295, 74.12193, 67.39835, 53.07862,
    56.73719, 57.33643, 59.6986, 62.59421, 65.6245, 66.04916, 65.75653,
    63.89017, 64.67288, 64.98264, 64.40124, 63.22442, 63.00884, 63.78863,
    62.93642, 61.06512, 57.83271, 61.37905, 68.36539, 62.30514, 42.51343,
    34.02612, 33.94305,
  71.61339, 71.45967, 70.79596, 69.67047, 72.01058, 66.07849, 60.36748,
    66.28746, 70.6358, 71.47134, 65.79163, 58.2507, 57.15454, 57.46554,
    57.18875, 57.88478, 58.51729, 58.51879, 58.81702, 60.6378, 64.28531,
    62.11525, 56.11677, 56.02638, 62.06122, 60.48186, 44.76373, 34.10906,
    34.59517, 33.88616,
  76.06219, 70.11452, 76.62918, 81.76781, 79.08326, 71.60304, 74.53799,
    68.53002, 62.74383, 62.07753, 57.0508, 54.21199, 55.91106, 55.81231,
    54.01177, 54.16204, 53.3418, 53.27484, 53.38055, 54.90707, 58.80135,
    58.52139, 55.28336, 60.7138, 63.06055, 50.56997, 34.67387, 36.43508,
    35.03525, 34.27125,
  105.0976, 109.2559, 112.8475, 113.5538, 111.8903, 104.5112, 80.72635,
    66.98259, 72.29562, 65.15216, 61.30484, 60.22741, 64.31725, 66.09761,
    60.97095, 51.44905, 52.53625, 52.50636, 52.89814, 55.01309, 58.39838,
    59.06407, 57.25477, 53.51372, 49.72158, 43.04906, 35.71508, 37.25259,
    36.19339, 35.05038,
  111.5573, 114.3369, 113.4627, 109.4496, 102.7618, 96.48325, 94.28093,
    93.05317, 82.82769, 83.28397, 87.39646, 84.48351, 82.65194, 82.00803,
    74.74152, 63.20746, 60.13597, 65.24895, 67.9061, 63.50343, 58.42068,
    53.33663, 48.13823, 42.02006, 38.23459, 37.15014, 35.96744, 35.46617,
    35.31631, 34.81673,
  106.9166, 98.12077, 92.90931, 87.30089, 84.85918, 87.57784, 92.67476,
    89.88757, 84.56673, 83.83954, 80.57889, 75.98874, 75.91945, 77.6424,
    76.54391, 74.52663, 69.60052, 66.24245, 64.25065, 58.54742, 48.80825,
    45.10094, 39.74097, 36.85263, 36.82729, 36.30761, 35.56477, 34.81523,
    34.43503, 34.15527,
  85.6012, 83.87698, 83.38844, 81.8982, 80.41156, 80.7343, 80.74597,
    76.97478, 72.50845, 68.70158, 66.86023, 64.821, 64.72071, 67.15653,
    64.646, 62.52252, 60.85892, 55.19759, 51.42986, 46.46376, 40.6752,
    39.65208, 37.06545, 36.41571, 36.61794, 36.24986, 35.47557, 34.91759,
    34.43684, 34.11047,
  75.27498, 73.73773, 72.61857, 71.50376, 70.14983, 68.36839, 67.11646,
    66.76243, 64.95029, 62.19457, 59.13473, 60.72354, 63.30431, 60.73591,
    56.16141, 53.41992, 50.74828, 48.07693, 46.76511, 44.12714, 39.50761,
    39.41971, 37.48134, 36.51226, 36.53061, 36.38536, 35.26591, 34.47638,
    34.18594, 34.04765,
  64.4977, 64.10291, 62.7787, 62.43514, 61.91817, 61.8145, 61.78158,
    62.35614, 62.55157, 61.06397, 62.07468, 63.26129, 61.58125, 59.44617,
    55.29262, 51.30793, 47.71462, 46.44462, 46.56284, 44.05408, 39.41459,
    39.02191, 37.60161, 36.78068, 36.12136, 35.78124, 35.11976, 34.201,
    33.99727, 33.91618,
  69.7717, 65.88938, 59.50148, 56.2317, 57.25999, 57.0579, 57.29113,
    57.53957, 56.84205, 56.92702, 58.02162, 56.04606, 51.75373, 50.96047,
    49.44036, 50.24975, 53.89998, 57.21555, 56.93913, 52.66301, 45.37854,
    40.98093, 38.56538, 37.70857, 36.5035, 35.86288, 35.21125, 34.29046,
    33.946, 33.9039,
  68.91637, 63.90494, 56.76474, 52.95063, 53.65168, 53.28047, 53.15342,
    53.03337, 53.47125, 55.18016, 54.87997, 51.32714, 50.84466, 50.13644,
    49.57591, 50.56773, 53.75139, 57.11436, 57.01944, 54.16719, 48.64818,
    43.5581, 40.29364, 39.14283, 37.82631, 36.47769, 35.52929, 34.46148,
    33.94825, 33.91718,
  66.35518, 61.96901, 54.60272, 50.92989, 51.44408, 51.28348, 51.37611,
    51.72644, 52.92439, 54.46885, 53.24413, 51.30712, 52.89547, 52.40854,
    51.24762, 50.6165, 50.64631, 50.61739, 49.93769, 47.67052, 45.90981,
    44.92451, 42.89281, 40.92834, 38.98108, 37.11015, 35.55653, 34.53058,
    33.99686, 33.93262,
  64.6172, 61.27254, 54.37671, 51.16132, 51.78517, 51.40576, 52.12075,
    52.84195, 54.47787, 54.80838, 52.11597, 50.49508, 50.9243, 50.03121,
    48.53816, 47.38474, 46.23644, 45.47788, 45.05844, 44.47661, 43.98273,
    43.45701, 43.39513, 42.40296, 40.243, 37.32102, 35.65573, 34.77179,
    34.12028, 33.97339,
  63.60529, 61.51311, 54.3806, 51.76118, 53.50658, 53.63063, 53.15228,
    52.18231, 52.27411, 50.78038, 47.56837, 47.01499, 46.81818, 46.30873,
    45.33951, 45.06444, 44.55456, 43.46692, 42.96165, 42.60984, 42.26204,
    41.70721, 41.19833, 41.14912, 41.01218, 38.32476, 36.12199, 35.45864,
    34.62933, 34.03122,
  65.58541, 64.63255, 59.79643, 57.88269, 57.90995, 56.55886, 56.15977,
    55.46544, 56.34565, 54.1575, 51.14768, 52.14025, 53.10177, 53.08815,
    51.73534, 50.78342, 49.46834, 47.51024, 45.67401, 44.52425, 43.65739,
    42.71952, 41.61409, 40.94692, 41.3423, 40.94509, 38.75026, 36.29799,
    35.42045, 34.43991,
  67.62704, 64.6883, 59.26537, 56.72518, 56.19182, 54.96385, 55.27212,
    57.70398, 60.92768, 58.67191, 55.60585, 56.93695, 57.91212, 58.10625,
    56.64405, 55.54456, 53.49121, 51.3777, 49.39441, 47.60583, 46.38915,
    44.69415, 42.5138, 41.29107, 41.6937, 42.24855, 41.39852, 38.22561,
    36.49454, 35.30468,
  68.89777, 66.73682, 61.72178, 57.81562, 56.50767, 55.79115, 58.31047,
    62.2846, 63.27495, 60.32929, 59.67392, 60.22634, 60.81031, 59.92587,
    57.79666, 56.50247, 54.85992, 52.96111, 51.16434, 49.3685, 48.11513,
    46.36716, 43.37612, 41.84997, 41.97508, 41.9312, 41.78939, 39.37185,
    36.3108, 35.13105,
  70.78951, 68.14038, 63.12216, 59.56196, 58.44668, 57.4946, 60.15317,
    62.23306, 61.82201, 60.14651, 60.50867, 60.76443, 60.93486, 60.04892,
    58.36575, 56.91676, 55.65952, 54.42358, 52.78905, 51.40545, 50.89089,
    50.33511, 48.28065, 46.0713, 45.14709, 44.55507, 44.3704, 41.97034,
    36.7971, 34.40841,
  71.79174, 69.30875, 65.55946, 64.2148, 65.01772, 64.40623, 63.97626,
    62.87634, 60.96881, 60.97907, 61.46361, 61.91224, 62.60023, 62.26752,
    60.84111, 59.17311, 57.77802, 56.83429, 56.13767, 55.29958, 53.64031,
    51.29649, 48.51261, 46.81405, 46.18111, 45.38503, 44.61273, 44.04791,
    40.64875, 35.32357,
  63.33677, 63.34274, 63.70261, 64.09788, 65.91952, 67.64297, 64.91557,
    59.91854, 58.39744, 58.53884, 58.07831, 57.93096, 57.97814, 57.87919,
    57.30699, 56.4643, 55.29744, 53.84334, 51.51336, 49.39819, 47.8182,
    46.235, 44.52732, 43.25908, 42.84577, 42.25583, 41.191, 39.72936,
    38.7129, 36.31305,
  57.99214, 58.52021, 58.81314, 58.59805, 60.3181, 63.48494, 63.10336,
    57.40504, 55.17607, 56.14127, 56.48248, 56.36833, 55.27987, 53.16432,
    51.07726, 49.58599, 46.84613, 44.54807, 43.43415, 42.0676, 40.94199,
    40.69325, 40.55083, 40.21022, 39.70744, 39.22124, 38.15678, 36.7103,
    35.47277, 34.23849,
  5.702757, 4.932442, 5.281432, 5.428281, 5.493974, 5.607255, 5.839027,
    6.149187, 6.650138, 7.605025, 9.356037, 11.36548, 12.69199, 15.81858,
    19.42963, 22.44545, 25.80302, 29.77943, 34.29395, 39.23032, 44.15641,
    48.1581, 51.12478, 53.0261, 53.90534, 53.89304, 53.56487, 54.4029,
    50.18037, 47.43177,
  5.046435, 4.565083, 4.748052, 5.33639, 5.605518, 5.78647, 6.161005, 6.3998,
    6.695465, 7.296906, 8.649919, 10.99585, 13.49228, 15.7306, 18.49722,
    21.87253, 25.7916, 30.24106, 35.09697, 40.45924, 45.27101, 49.40108,
    52.39608, 54.29311, 55.03525, 54.42293, 53.14177, 54.13233, 50.29045,
    48.10794,
  7.765629, 7.82601, 8.776732, 9.399588, 9.943777, 10.05947, 10.16135,
    10.26763, 10.43006, 10.77428, 11.48269, 12.6828, 14.49163, 16.91839,
    19.69707, 22.80156, 26.551, 31.0989, 36.27254, 41.89103, 47.22624,
    51.6605, 54.66954, 55.98405, 56.02361, 55.48433, 54.97255, 53.93917,
    49.40343, 47.97613,
  10.36386, 9.542824, 9.900473, 9.889318, 10.0235, 10.18069, 10.30332,
    10.43322, 10.75788, 11.36186, 12.3602, 13.63743, 15.31928, 17.68414,
    20.59401, 23.76469, 27.30124, 31.23215, 36.39106, 41.98616, 47.47746,
    51.82044, 54.35907, 56.16671, 56.3912, 56.46053, 56.42847, 55.29255,
    53.90878, 48.60899,
  10.83444, 10.04062, 10.43895, 10.40282, 10.44119, 10.43486, 10.48849,
    10.54732, 10.88505, 11.66199, 12.92391, 14.68168, 16.68261, 19.07399,
    21.91807, 25.15146, 28.74481, 32.70035, 37.49132, 43.08282, 47.85185,
    51.22058, 53.96798, 55.56591, 56.0764, 56.10613, 56.00326, 56.87426,
    56.40055, 54.22409,
  10.67745, 10.15781, 10.69793, 10.9211, 10.98565, 10.94804, 11.16628,
    11.32497, 11.38661, 11.78705, 12.86036, 14.62897, 17.18263, 19.69409,
    22.64602, 26.19158, 30.39705, 34.67072, 39.20786, 44.37364, 48.5697,
    51.62277, 54.24387, 55.39828, 55.66473, 55.47829, 55.1571, 55.74304,
    55.66299, 52.50722,
  10.67145, 10.07281, 10.63558, 10.89114, 11.16147, 11.4057, 11.77589,
    12.21757, 12.59301, 12.992, 13.7232, 14.61494, 15.73891, 18.28652,
    21.36466, 25.01411, 29.22072, 34.02779, 38.73785, 44.24142, 48.80812,
    52.23745, 54.57455, 55.80904, 55.92407, 55.33736, 55.15246, 55.29658,
    54.58352, 45.77753,
  11.50734, 10.52269, 10.98184, 11.07616, 11.22396, 11.66562, 12.03149,
    11.1241, 10.93599, 11.80654, 12.90478, 14.42976, 16.40088, 18.90115,
    21.92912, 25.19293, 29.39728, 34.26071, 39.15398, 44.28352, 49.01878,
    52.63948, 54.93064, 55.93589, 55.77984, 55.56654, 55.72062, 55.26165,
    53.84231, 46.16156,
  14.59218, 12.77209, 12.55069, 12.23343, 12.01044, 11.89544, 10.92078,
    10.86668, 11.1938, 11.93939, 13.28962, 15.04254, 17.05487, 19.76571,
    22.98737, 25.61342, 29.63084, 34.90316, 40.28476, 45.19948, 49.55678,
    53.14746, 55.21891, 55.69777, 55.37265, 55.75945, 55.77273, 54.70848,
    46.6663, 46.87518,
  19.95448, 17.8445, 16.37622, 15.18966, 14.55762, 13.4674, 11.48351,
    11.7281, 11.71017, 12.25755, 13.56509, 15.96467, 18.21441, 19.97265,
    22.41187, 26.05201, 30.13363, 34.79344, 39.9289, 45.36073, 50.32771,
    53.48092, 54.64438, 54.44201, 54.78555, 55.26212, 54.97947, 53.33524,
    46.08127, 45.73242,
  24.93979, 22.42983, 22.32689, 20.00158, 18.76994, 16.75719, 14.92205,
    13.685, 13.36218, 14.08906, 14.67151, 16.16648, 17.77143, 20.05219,
    22.89029, 26.03039, 29.93895, 34.40244, 39.30463, 44.41085, 50.01845,
    53.39111, 54.33003, 54.37937, 54.78486, 54.52182, 53.34617, 46.76816,
    47.16781, 45.83736,
  24.96332, 22.88401, 25.65472, 26.07581, 24.93381, 21.29149, 17.97649,
    14.70525, 13.235, 13.82837, 14.82472, 16.45123, 19.00179, 21.07568,
    23.37642, 26.85281, 30.24886, 34.70626, 39.58715, 44.43539, 49.33012,
    53.07587, 54.05211, 54.73897, 55.02431, 54.18524, 46.91246, 51.58788,
    47.98426, 46.62199,
  14.84516, 16.31137, 18.68671, 21.71193, 24.01231, 23.67094, 17.32746,
    12.04876, 15.72902, 14.41626, 15.79606, 16.87544, 18.98319, 21.33824,
    24.02395, 26.49402, 30.60678, 35.12648, 40.00507, 45.02367, 49.56821,
    52.56946, 53.87394, 53.72902, 53.71918, 53.40633, 47.69884, 49.35464,
    48.88768, 47.47814,
  11.3238, 10.06414, 10.17167, 10.40825, 10.97941, 11.84328, 12.86821,
    14.07503, 12.99842, 14.12545, 15.88648, 17.79673, 19.59816, 21.63586,
    24.45754, 27.2191, 30.3194, 35.60664, 40.90567, 45.5885, 49.11325,
    51.91655, 53.08941, 50.61933, 47.2784, 47.59194, 46.97701, 46.50019,
    46.78262, 46.80005,
  12.26285, 11.17006, 11.67461, 11.71123, 11.96891, 12.09256, 12.38673,
    12.51227, 12.90889, 14.11496, 15.7486, 17.64949, 19.76449, 22.12681,
    24.18809, 26.91366, 30.8249, 34.1658, 39.74672, 45.0563, 48.28258,
    51.22057, 50.6767, 48.56374, 48.87634, 48.02275, 47.21594, 46.66264,
    46.11884, 45.95802,
  10.92295, 10.53229, 11.05381, 11.2994, 11.73439, 12.30653, 12.99591,
    13.24122, 13.70993, 15.21408, 17.36694, 19.22863, 21.19644, 22.85547,
    24.90158, 27.53986, 30.45774, 33.94957, 39.24861, 44.4531, 45.85498,
    49.19037, 48.96471, 48.75619, 48.5626, 47.86164, 47.05811, 46.62807,
    46.18912, 45.98495,
  8.046144, 6.445599, 8.097462, 9.788727, 10.58551, 11.08275, 11.67362,
    12.39908, 13.52677, 15.26459, 17.29289, 20.01568, 23.12885, 25.13466,
    27.30734, 29.50243, 31.96198, 35.55816, 40.79161, 45.22512, 46.20358,
    49.37971, 49.19189, 48.75932, 48.64916, 48.13442, 47.02256, 46.10925,
    45.86002, 45.8752,
  11.42142, 8.249321, 7.028687, 7.40904, 8.653678, 9.841996, 10.65232,
    11.10276, 11.93633, 13.19136, 15.65039, 18.75556, 21.6785, 25.74291,
    29.07232, 31.67997, 34.47095, 38.57036, 43.62787, 47.79824, 49.39038,
    49.70668, 49.38377, 49.23389, 48.52144, 47.99656, 47.24725, 46.06425,
    45.70752, 45.72518,
  22.00889, 16.93906, 10.23972, 4.85024, 6.942721, 7.0845, 8.079359,
    9.128966, 10.18741, 12.18995, 14.28305, 16.47178, 19.00169, 22.71017,
    27.27795, 31.18825, 35.67033, 41.31274, 47.30702, 51.69178, 53.56598,
    53.91402, 51.10096, 50.78413, 49.38671, 48.45102, 47.59126, 46.27605,
    45.66478, 45.76208,
  21.44928, 16.91935, 10.44703, 5.40626, 6.906943, 7.207491, 8.183736,
    9.300018, 11.07516, 12.89865, 14.42833, 15.68651, 18.2498, 20.88577,
    24.15356, 28.54816, 33.39769, 39.02021, 45.17765, 50.18269, 53.65497,
    55.05089, 53.42545, 52.19844, 50.60222, 48.98799, 47.79414, 46.40764,
    45.64895, 45.77955,
  22.26883, 17.78965, 12.39043, 7.604733, 8.611301, 8.619959, 9.488789,
    10.52618, 12.25106, 13.72043, 14.58857, 15.264, 19.11197, 21.73541,
    24.59983, 28.20484, 33.12916, 38.52419, 43.92951, 48.74451, 52.37468,
    54.8496, 55.68547, 54.0127, 51.8762, 49.59416, 47.85425, 46.41621,
    45.67459, 45.78788,
  23.13435, 19.34649, 14.96629, 12.29705, 13.46284, 13.25448, 13.83777,
    14.1608, 14.96523, 15.9684, 16.81074, 17.76661, 20.97769, 23.78769,
    26.66251, 30.33724, 34.50209, 39.48185, 44.32162, 48.62809, 52.2595,
    54.60228, 55.79038, 55.8268, 54.1002, 50.6705, 48.4093, 46.95966,
    45.84232, 45.78792,
  23.3368, 20.08628, 16.18703, 14.05751, 15.56199, 16.0999, 16.78812,
    17.32815, 18.31147, 19.39154, 20.70371, 22.93602, 25.45224, 28.0493,
    30.79846, 34.1715, 38.14756, 42.38174, 46.63912, 50.38959, 53.35559,
    55.05917, 55.45265, 55.76411, 55.81446, 53.09323, 49.75332, 47.99611,
    46.70352, 45.93912,
  23.27962, 19.91868, 16.54323, 14.90235, 16.15645, 16.76551, 18.09026,
    19.60361, 21.33186, 22.44772, 24.2522, 27.47188, 31.15465, 34.27498,
    36.76402, 39.81822, 43.24149, 46.91492, 50.60133, 54.02338, 56.38021,
    57.41462, 56.91374, 56.43253, 56.6884, 56.07204, 53.33571, 49.61581,
    48.08714, 46.74869,
  23.05028, 19.09129, 15.47039, 13.39763, 14.56247, 15.2083, 16.6325,
    18.59487, 20.53876, 21.74227, 23.42905, 26.83871, 30.79628, 34.21717,
    36.71648, 39.99218, 43.47163, 47.25282, 51.21914, 54.98319, 57.52322,
    58.53219, 57.91927, 56.28224, 56.40692, 56.27866, 55.08304, 51.42813,
    48.82063, 47.62349,
  24.99584, 21.04809, 17.30547, 15.02097, 15.76002, 16.25247, 17.7626,
    19.76209, 21.41903, 22.70474, 24.85656, 28.0253, 31.80821, 34.80652,
    37.08272, 40.09887, 43.38029, 47.00739, 50.97827, 54.81952, 57.59261,
    58.92588, 58.3746, 57.57681, 57.29434, 56.53706, 55.49418, 52.33634,
    48.36095, 47.07319,
  32.37145, 28.79617, 25.01173, 22.7784, 23.53272, 23.69962, 24.99515,
    26.42213, 27.64609, 28.87427, 31.00199, 33.81964, 37.20366, 39.81565,
    41.55357, 43.68773, 46.00452, 48.84496, 52.13709, 55.41659, 57.8232,
    59.05839, 58.89999, 58.1293, 57.77121, 57.1224, 56.33455, 54.8645,
    50.12828, 46.71021,
  42.99171, 41.26569, 38.33, 36.88837, 37.77717, 38.03594, 38.6215, 39.2578,
    39.64684, 40.22409, 41.19318, 42.75693, 45.11421, 47.00952, 47.93846,
    49.11362, 50.26268, 51.62632, 53.72564, 56.048, 57.57053, 58.19323,
    57.15395, 56.25121, 56.3712, 56.05614, 55.4591, 54.83302, 53.0412, 48.1717,
  46.99296, 47.29128, 47.52036, 48.21885, 49.01604, 49.85929, 50.00617,
    49.38499, 48.0313, 48.42414, 48.20018, 48.38881, 48.95626, 49.58131,
    49.85743, 50.10581, 50.07985, 50.26631, 50.50194, 51.09017, 51.92423,
    52.78004, 52.85722, 51.95434, 52.13371, 52.25146, 51.6362, 49.92671,
    49.2541, 48.21242,
  50.7961, 51.44374, 51.80414, 51.89585, 53.07767, 53.99894, 54.56449,
    52.29597, 49.94173, 50.73974, 51.16897, 51.92496, 51.9649, 51.42958,
    50.61586, 50.09925, 48.9759, 47.64158, 47.54205, 47.71976, 47.58311,
    48.32807, 49.16269, 49.52214, 49.60321, 49.86893, 49.51831, 48.16754,
    46.9521, 46.00493,
  22.02957, 23.8093, 25.99256, 28.22123, 30.67991, 33.19903, 35.88983,
    38.59977, 41.45059, 44.36954, 47.27533, 49.85342, 51.75676, 53.23397,
    54.23803, 54.90474, 55.3063, 55.58124, 55.84869, 56.21543, 56.46345,
    56.42039, 56.38581, 56.37894, 56.11528, 55.37306, 51.96374, 55.24892,
    50.97, 47.77236,
  21.23301, 23.05568, 25.47121, 27.95508, 30.44428, 33.22021, 36.21209,
    39.21108, 42.14794, 45.08722, 48.05005, 50.73259, 52.8888, 54.21708,
    54.90854, 55.37098, 55.50924, 55.68698, 55.97574, 56.47939, 57.04334,
    57.57383, 57.87489, 58.04232, 58.00211, 56.87872, 55.17216, 53.31765,
    50.11955, 48.03796,
  21.91776, 23.73995, 26.12752, 28.58979, 30.93568, 33.66328, 36.67877,
    39.8531, 42.94092, 45.84348, 48.57453, 51.14817, 53.32648, 54.82992,
    55.67433, 55.85561, 55.83735, 55.90742, 56.00994, 56.28419, 57.02296,
    57.9123, 58.38498, 58.55945, 58.29792, 58.08062, 57.41061, 55.59455,
    50.57579, 47.64926,
  22.35229, 24.22553, 27.14776, 29.40822, 31.8097, 34.19865, 36.8562,
    39.93994, 43.16975, 46.32395, 49.15757, 51.68756, 53.90392, 55.36587,
    56.24343, 56.57019, 56.44755, 56.2578, 56.46715, 56.73951, 57.21095,
    57.35139, 56.94289, 57.58327, 57.59389, 58.06401, 58.41485, 57.69208,
    55.86029, 50.81325,
  23.08152, 24.84605, 27.5943, 30.38522, 32.75795, 35.04503, 37.30579,
    40.17111, 43.0111, 46.13626, 49.14489, 51.89725, 54.42013, 56.05846,
    57.00934, 57.36385, 57.18887, 56.8949, 56.95461, 57.2933, 57.15542,
    56.42585, 56.6555, 57.03191, 57.25631, 57.39489, 57.57452, 58.70089,
    58.34944, 55.8052,
  24.31342, 25.60671, 28.21252, 30.8604, 33.60794, 35.93637, 38.07654,
    41.12957, 43.72498, 46.19672, 48.88257, 51.66711, 54.46111, 56.15321,
    57.30448, 57.96299, 57.75442, 57.45998, 57.1301, 57.16468, 56.81702,
    56.09745, 56.84881, 57.2259, 57.24829, 57.17096, 57.00354, 57.59658,
    57.51424, 53.19316,
  27.68298, 27.85654, 29.51015, 31.53274, 33.97234, 36.54678, 38.83719,
    41.71983, 44.69252, 47.12769, 49.45659, 51.31796, 52.49693, 54.33204,
    55.53062, 56.29097, 56.72731, 56.53483, 55.9074, 55.95124, 56.02919,
    56.20903, 56.70678, 57.31055, 57.44008, 57.26044, 57.34963, 57.36315,
    56.39671, 45.97406,
  33.2815, 32.52557, 32.88082, 33.69253, 35.27851, 37.79223, 40.20545,
    41.22701, 43.17141, 45.75731, 48.07283, 50.23905, 52.26315, 54.16796,
    55.52518, 56.23231, 56.89016, 57.17123, 56.77745, 56.26269, 56.07317,
    56.29531, 56.67612, 57.01633, 57.09933, 57.36276, 57.65046, 56.9448,
    55.20055, 46.35433,
  38.98635, 39.29536, 38.67654, 38.37791, 38.7344, 39.79703, 40.05383,
    42.09236, 44.58531, 46.78541, 48.84187, 50.71083, 52.26294, 53.96378,
    55.54644, 56.02441, 56.67255, 57.43147, 57.84348, 57.34749, 56.78658,
    56.55333, 56.61092, 56.45444, 56.42946, 57.1307, 57.36718, 56.21625,
    46.23518, 46.9615,
  41.16522, 44.29845, 45.20721, 44.73345, 43.93225, 43.19829, 42.00073,
    43.62471, 45.58961, 47.9457, 49.63959, 51.45932, 52.69368, 53.57135,
    54.32983, 55.35559, 56.00762, 56.59173, 57.04773, 57.20351, 57.40923,
    56.78265, 56.29293, 55.77932, 56.15788, 56.56456, 56.37188, 54.17221,
    46.50679, 46.09981,
  38.87351, 42.10661, 46.96122, 49.31752, 49.62383, 47.82215, 46.51455,
    46.23251, 46.78328, 49.39731, 50.73669, 51.6908, 52.67, 53.47675,
    54.11673, 54.78436, 55.27368, 55.69225, 56.1323, 56.37658, 57.0667,
    56.73815, 55.92492, 56.04768, 56.73742, 56.35471, 54.68851, 48.46321,
    47.82385, 46.41251,
  34.94371, 34.87222, 42.0698, 47.93974, 52.97546, 52.04905, 49.22131,
    46.97227, 48.0178, 49.36875, 51.22489, 52.47114, 54.03893, 54.73682,
    54.82375, 54.9731, 55.53239, 55.94213, 56.14323, 56.14737, 56.71303,
    56.69508, 55.61086, 55.71997, 56.47574, 55.98432, 46.70611, 53.40214,
    49.0449, 47.38134,
  29.2274, 31.5374, 34.11166, 39.58126, 45.95932, 50.76982, 48.44186,
    45.03982, 50.70472, 51.04494, 52.96721, 54.0428, 55.43282, 56.45552,
    56.53983, 55.20861, 55.74366, 56.4648, 56.72017, 56.39293, 56.54534,
    56.43835, 55.71732, 54.83841, 54.81838, 54.80881, 47.64536, 49.0019,
    49.57722, 48.20801,
  27.81875, 29.52141, 31.0315, 33.25599, 35.75214, 38.81149, 43.2336,
    47.70163, 48.59196, 51.24815, 53.74906, 55.71499, 56.62115, 57.44309,
    57.54198, 56.60032, 55.85065, 56.47151, 57.15996, 56.52342, 55.66564,
    55.42082, 54.80708, 51.42558, 47.09299, 47.51827, 47.56586, 46.55003,
    46.87618, 47.30802,
  26.05137, 27.14423, 30.32868, 33.28439, 36.22455, 39.10536, 41.65901,
    44.6068, 48.12553, 50.93219, 53.10448, 54.92179, 56.59519, 57.82911,
    58.05413, 58.06599, 57.1763, 56.04363, 55.67513, 55.53191, 54.46395,
    54.51717, 51.73351, 48.72923, 49.23521, 48.26205, 47.65607, 47.17773,
    46.46831, 46.3097,
  25.2221, 27.40517, 29.41851, 31.57021, 34.38813, 37.26296, 40.27509,
    43.26181, 46.39364, 49.7264, 52.4177, 54.54413, 56.45837, 58.14219,
    58.76383, 58.689, 58.44943, 57.28173, 56.1075, 55.28458, 52.73379,
    52.59978, 50.43984, 49.14043, 48.82517, 48.15426, 47.2988, 46.88316,
    46.50891, 46.37351,
  28.34892, 27.68701, 30.55043, 32.58926, 34.90074, 37.48078, 40.13957,
    42.43506, 45.21402, 48.16637, 50.78099, 53.58865, 56.1723, 57.70927,
    58.76443, 59.5692, 59.93737, 59.77362, 58.68545, 57.0815, 54.70544,
    53.30191, 51.2247, 49.77197, 49.32839, 48.71342, 47.42361, 46.40404,
    46.20436, 46.22572,
  35.58883, 33.00045, 32.92517, 33.93727, 36.88338, 39.01827, 41.61544,
    44.01607, 46.02618, 48.33278, 50.90341, 53.33159, 54.92392, 56.43076,
    57.45925, 58.61162, 59.9501, 61.07241, 61.47295, 60.25768, 57.6235,
    55.34917, 52.283, 51.08279, 49.59976, 48.90979, 47.85136, 46.47512,
    46.15126, 46.11916,
  46.16431, 41.76067, 37.62803, 35.16841, 38.71188, 40.91497, 43.44831,
    45.9015, 48.54532, 50.69074, 52.85605, 54.45578, 55.35064, 55.9787,
    56.28931, 56.93664, 58.31639, 60.0867, 61.23684, 61.60466, 60.51102,
    58.12434, 54.77092, 53.44678, 51.01041, 49.77837, 48.5249, 46.82483,
    46.11226, 46.1552,
  45.8716, 42.67268, 38.60429, 36.85238, 40.15054, 42.3218, 45.29334,
    47.98557, 50.67812, 53.04836, 54.99498, 56.25969, 57.58769, 57.98478,
    57.88297, 57.69438, 57.84578, 58.4034, 58.72926, 58.95797, 59.38762,
    58.84229, 57.37878, 55.15739, 52.85888, 50.56904, 48.99135, 47.02048,
    46.04953, 46.16786,
  47.66939, 44.0677, 40.1871, 38.791, 42.18399, 44.40129, 47.3171, 50.33205,
    53.19963, 55.69967, 57.43335, 58.60655, 59.90272, 60.53302, 60.39137,
    60.09776, 59.82371, 59.7098, 59.318, 58.54635, 58.36681, 58.57149,
    58.26144, 57.24656, 54.7574, 51.71968, 49.29018, 47.28651, 46.02525,
    46.14166,
  50.59213, 47.53004, 43.18958, 41.58535, 45.24546, 47.46315, 50.33595,
    53.0041, 56.01727, 58.76473, 60.84338, 62.38841, 63.41547, 63.90815,
    63.71375, 63.04079, 62.21317, 61.56911, 60.82206, 59.80056, 59.35057,
    58.82251, 58.77381, 58.15675, 57.06424, 53.56901, 50.17405, 48.16418,
    46.44299, 46.11467,
  55.93907, 52.61161, 48.33183, 46.4243, 49.474, 51.74664, 54.49825,
    56.96639, 59.53064, 61.92385, 64.29061, 66.84763, 68.51817, 69.0983,
    68.70131, 67.96761, 66.70344, 65.25879, 63.80152, 62.42871, 61.37934,
    60.52785, 59.66428, 58.92324, 58.39108, 56.23542, 52.12275, 49.4437,
    47.67914, 46.46718,
  62.73611, 59.05791, 54.22393, 51.9849, 54.08205, 55.38073, 57.82248,
    60.52478, 63.38787, 65.0504, 66.87717, 70.03265, 73.29208, 74.38513,
    73.73209, 73.18971, 72.02802, 70.16669, 67.97729, 66.37922, 65.03792,
    63.39751, 61.33543, 60.15418, 59.80296, 58.74667, 55.76371, 51.01236,
    49.12237, 47.4892,
  68.14692, 63.46755, 58.18847, 55.11734, 56.31207, 56.7923, 58.41189,
    60.92788, 63.70134, 64.8958, 66.28591, 69.10671, 72.18776, 73.41649,
    72.42395, 72.40271, 71.66045, 70.42937, 68.69601, 67.23405, 66.07285,
    64.46829, 61.9591, 60.47506, 60.23823, 59.3685, 57.17036, 52.74662,
    49.3187, 48.16068,
  70.54475, 65.75792, 60.19682, 57.02886, 57.55802, 57.40427, 58.61161,
    60.55796, 62.27472, 62.84068, 64.42717, 67.32011, 70.40009, 71.19992,
    70.21324, 70.09191, 69.69753, 68.75631, 67.71416, 66.85089, 65.72641,
    64.30701, 62.04372, 60.5517, 60.34278, 59.46112, 58.12659, 54.1687,
    49.33371, 47.64346,
  69.42403, 65.55561, 60.43683, 57.39571, 58.03687, 57.73849, 58.47366,
    59.48558, 60.15905, 60.05564, 61.08426, 63.2403, 66.47492, 67.82294,
    67.08392, 66.84734, 66.32452, 65.92736, 65.54731, 65.34702, 64.7511,
    63.61441, 61.85758, 60.22234, 59.80169, 59.1537, 58.24942, 56.39777,
    51.25836, 47.63033,
  63.75787, 62.11029, 58.77024, 56.69444, 57.51333, 57.67799, 58.17403,
    58.59306, 57.67018, 57.38976, 57.15245, 58.59076, 60.63265, 62.23341,
    62.08849, 61.9375, 61.86835, 60.8229, 60.82083, 61.70113, 61.72261,
    60.55373, 58.03094, 56.38493, 56.23703, 55.54465, 54.54171, 53.63604,
    52.33646, 48.61731,
  53.25842, 54.08787, 54.76873, 55.12683, 55.62139, 56.2879, 56.60025,
    54.22533, 53.09904, 53.60858, 53.05458, 52.55028, 52.37902, 52.97876,
    53.16104, 53.08033, 52.4068, 51.69057, 50.98222, 50.8374, 51.50743,
    52.39633, 52.806, 52.12813, 52.51385, 52.59529, 51.75672, 49.7566,
    48.58524, 48.09078,
  50.23841, 50.52779, 50.95726, 51.0126, 51.79148, 53.48025, 54.21831,
    51.66801, 49.75528, 50.402, 50.752, 50.94687, 50.58064, 50.36272,
    50.08873, 49.89973, 48.94083, 47.62158, 47.45203, 47.45504, 47.15624,
    47.66791, 48.57155, 49.11948, 49.25251, 49.58033, 49.38581, 48.25126,
    47.07619, 46.35728,
  51.50694, 52.80258, 53.72439, 54.54108, 55.05418, 55.45626, 55.75187,
    55.92556, 56.03561, 56.19421, 56.37354, 56.51871, 56.56894, 56.79992,
    57.02457, 57.41046, 57.93325, 58.54156, 59.37244, 60.21652, 61.06221,
    61.57539, 61.86247, 62.07347, 61.86553, 56.09586, 51.08371, 53.53575,
    50.71138, 48.47361,
  51.19072, 52.49942, 53.43434, 54.3627, 54.9395, 55.36757, 55.69082,
    55.93204, 56.1451, 56.29441, 56.45466, 56.72026, 56.98407, 57.11525,
    57.10994, 57.38214, 57.75715, 58.36084, 59.25436, 60.40502, 61.6218,
    62.65963, 63.36474, 63.61264, 63.39657, 61.95578, 53.90033, 51.50193,
    50.12405, 48.69838,
  51.39731, 52.61898, 53.48816, 54.40332, 55.05534, 55.51152, 55.76827,
    56.04844, 56.33091, 56.52758, 56.72992, 57.04152, 57.34803, 57.59655,
    57.80175, 57.87783, 58.09242, 58.51525, 59.17736, 60.14131, 61.52992,
    63.04557, 63.9162, 64.23512, 63.90709, 63.03681, 62.11998, 57.27192,
    50.04392, 48.60736,
  51.58004, 52.68059, 53.54395, 54.40709, 55.10108, 55.6941, 55.99839,
    56.16391, 56.38023, 56.61512, 56.96199, 57.49585, 57.85239, 57.99286,
    58.31603, 58.61548, 58.73574, 58.95181, 59.57104, 60.4137, 61.48703,
    62.30024, 62.47851, 63.27985, 63.34134, 63.63228, 63.4377, 62.7086,
    61.45818, 50.9025,
  51.83604, 52.87965, 53.75961, 54.5099, 55.08717, 55.72229, 56.27692,
    56.42418, 56.42662, 56.54827, 57.06441, 57.93116, 58.57879, 58.7733,
    59.05723, 59.44174, 59.59309, 59.63486, 60.14426, 60.83778, 61.20029,
    61.22914, 61.96095, 62.73995, 63.12234, 63.08577, 63.21949, 64.14971,
    63.87042, 61.7486,
  52.50712, 53.26078, 54.21169, 54.86426, 55.23977, 55.73132, 56.48595,
    56.92538, 56.97063, 56.98895, 57.35771, 58.09647, 58.99578, 59.14264,
    59.52058, 59.98874, 59.97102, 60.12464, 60.44672, 60.80563, 60.88409,
    60.73463, 61.96147, 62.66216, 62.87455, 62.81644, 62.70887, 63.15228,
    63.07667, 53.73547,
  54.57756, 54.2806, 54.95222, 55.38713, 55.68288, 56.0733, 56.69342,
    56.93526, 57.19559, 57.42606, 57.69759, 57.53087, 56.93497, 57.51458,
    57.98679, 58.37245, 58.72172, 58.93011, 59.09594, 59.6647, 60.08401,
    60.75322, 61.7668, 62.67384, 62.9891, 62.90678, 63.01609, 63.05949,
    62.12803, 47.29595,
  58.91539, 57.30584, 56.85333, 56.70674, 56.67668, 56.94065, 57.16677,
    56.02991, 55.40578, 55.61796, 55.87921, 56.21117, 56.69514, 57.38338,
    58.01639, 58.48577, 58.99754, 59.46843, 59.64596, 59.75126, 60.07368,
    60.79666, 61.71524, 62.43081, 62.66002, 63.0353, 63.24377, 62.60183,
    61.20213, 47.60652,
  64.48443, 63.16342, 61.11971, 59.73672, 58.68151, 57.965, 56.46597,
    56.52118, 56.41548, 56.03477, 56.03391, 56.27412, 56.50328, 57.18959,
    58.01179, 58.38379, 59.13195, 60.10228, 60.79886, 60.7077, 60.72906,
    61.09334, 61.63136, 61.89251, 62.09174, 62.80372, 63.09303, 61.94466,
    47.57065, 48.16459,
  67.23475, 68.74941, 67.32741, 65.22351, 63.05822, 60.4044, 57.67128,
    57.53568, 57.26988, 57.09886, 56.60676, 56.58344, 56.60233, 56.75627,
    57.07237, 57.84661, 58.63697, 59.55783, 60.40921, 60.87192, 61.33069,
    61.35423, 61.39186, 61.47097, 62.01659, 62.2413, 61.95469, 54.39266,
    47.57197, 47.59264,
  64.89536, 67.65987, 70.87931, 70.70233, 69.01441, 64.74192, 61.43272,
    59.22783, 58.0934, 58.52714, 57.59739, 56.76108, 56.61555, 56.68818,
    56.90721, 57.44035, 58.06466, 58.79911, 59.61448, 60.2719, 61.13171,
    61.40555, 61.39825, 61.93665, 62.91519, 62.63271, 57.20933, 48.65338,
    48.75249, 47.75633,
  60.60364, 60.7401, 66.23589, 70.33508, 71.867, 68.72723, 64.28105,
    60.52053, 59.05941, 58.85805, 58.33032, 57.80197, 57.95736, 57.81087,
    57.39209, 57.56269, 58.23221, 58.944, 59.54185, 60.03111, 60.83499,
    61.28776, 61.18403, 61.74112, 62.59049, 62.15986, 48.10717, 53.62448,
    49.66405, 48.431,
  54.76064, 56.40518, 58.16313, 61.52307, 65.13271, 66.77351, 62.26493,
    58.64746, 61.35789, 60.1389, 59.79178, 59.12715, 59.29928, 59.40961,
    58.8618, 57.65395, 58.4222, 59.37131, 59.98926, 60.24869, 60.9378,
    61.35547, 61.22609, 57.90141, 56.61532, 58.08503, 48.62324, 50.20776,
    50.34051, 49.17164,
  55.13923, 55.63241, 55.63374, 55.17237, 55.23414, 56.54383, 58.6773,
    60.19225, 58.87777, 59.89952, 60.48902, 60.22953, 60.03629, 60.09376,
    59.5206, 58.50443, 58.23184, 59.21678, 60.30083, 60.44379, 60.5004,
    60.73812, 56.12909, 51.43646, 47.93111, 48.55888, 48.57012, 47.80989,
    48.20401, 48.5112,
  55.42848, 55.97472, 56.60187, 56.74262, 56.956, 57.33681, 57.87797,
    58.0524, 58.28288, 58.58152, 59.04647, 59.3449, 59.77735, 60.04398,
    59.76659, 59.49495, 58.8578, 58.51289, 58.8875, 59.42356, 55.76169,
    55.54241, 52.05795, 49.08913, 49.82148, 49.28482, 48.78703, 48.29593,
    47.81277, 47.71465,
  56.01122, 56.62321, 57.05965, 57.05317, 57.08185, 57.59716, 58.09817,
    58.19651, 57.97433, 58.06349, 58.58204, 59.25945, 60.01459, 60.75319,
    60.59283, 60.05309, 59.91781, 59.3962, 56.92122, 54.95206, 52.90207,
    52.29987, 50.46171, 49.39321, 49.31177, 49.02696, 48.50124, 48.22287,
    47.89322, 47.8346,
  58.37322, 58.12865, 58.44526, 58.58892, 58.50642, 58.29654, 58.34996,
    58.55301, 58.34185, 58.04944, 58.03939, 58.86351, 60.10112, 60.87895,
    61.29993, 61.6091, 61.85946, 61.8527, 61.13488, 58.56496, 53.79758,
    52.8725, 51.30885, 50.1229, 49.92597, 49.40478, 48.50478, 47.84095,
    47.67249, 47.69154,
  64.51611, 62.12767, 60.48015, 60.04766, 60.39808, 60.1042, 59.93711,
    59.6779, 59.46346, 58.8974, 58.77039, 58.90966, 59.09648, 59.67068,
    60.34681, 61.37524, 62.71481, 63.77186, 63.9109, 62.84376, 58.89967,
    54.22446, 52.33869, 51.52631, 50.63085, 49.95025, 48.85463, 47.86197,
    47.62482, 47.60451,
  74.02455, 69.42108, 64.26308, 60.88454, 62.25798, 61.82932, 61.71535,
    61.36502, 60.7245, 60.44773, 60.34927, 60.05534, 59.47366, 58.84507,
    58.30115, 59.66245, 61.19946, 63.1025, 64.38525, 64.82848, 63.98616,
    58.99416, 54.26712, 53.68036, 51.89558, 50.82829, 49.67395, 48.22583,
    47.58251, 47.63271,
  73.63772, 69.67516, 64.41277, 62.01426, 63.2483, 63.2832, 63.31671,
    62.99532, 62.5101, 62.04717, 61.79921, 61.52523, 61.40951, 60.70837,
    59.85685, 58.42212, 58.49809, 60.4268, 62.04634, 62.70697, 63.2317,
    61.09806, 56.7179, 54.82747, 53.16681, 51.35612, 50.06576, 48.39735,
    47.54563, 47.64087,
  73.82257, 70.11908, 64.85265, 62.41225, 63.89439, 64.17885, 64.67997,
    64.81288, 64.74928, 64.28281, 63.70309, 63.06345, 62.85213, 62.5744,
    62.10102, 61.832, 61.8811, 62.14473, 61.81329, 60.19017, 59.31487,
    59.76978, 58.7789, 56.35396, 54.55828, 52.09035, 50.20227, 48.52306,
    47.48233, 47.58346,
  72.50637, 69.95355, 64.32346, 62.04894, 63.89179, 64.51217, 65.45774,
    66.0735, 66.68674, 67.02039, 66.64546, 65.9611, 65.2822, 64.70139,
    64.33355, 64.02837, 63.78013, 63.87699, 63.85099, 61.66408, 59.6459,
    58.33547, 59.18592, 57.62753, 56.35406, 53.64792, 51.02298, 49.0787,
    47.71431, 47.54705,
  71.0906, 68.47021, 63.46938, 60.83168, 62.93856, 64.01728, 65.3743,
    66.4215, 67.81838, 68.81846, 69.4249, 69.92622, 69.70409, 69.18803,
    68.44102, 67.94908, 67.45372, 67.0022, 66.42104, 65.5257, 62.79835,
    60.71328, 59.61208, 58.276, 58.16406, 56.13397, 52.9255, 50.23405,
    48.66563, 47.77776,
  70.87981, 67.29063, 62.11765, 59.80253, 61.26706, 62.327, 64.05284,
    66.17088, 68.42539, 69.45911, 70.54784, 72.11859, 74.33658, 74.61205,
    73.75074, 73.28949, 72.54465, 71.46613, 70.17621, 69.0348, 68.2472,
    65.80726, 62.17785, 60.22115, 59.99173, 59.05098, 56.27254, 51.93731,
    50.00157, 48.66666,
  70.95628, 66.44543, 61.43198, 58.49355, 59.30175, 59.89437, 61.71918,
    64.27498, 67.05174, 67.90594, 68.77567, 70.52693, 72.62939, 74.22649,
    73.58817, 73.61136, 73.23776, 72.32186, 71.01968, 70.28092, 69.39114,
    67.31784, 63.39039, 60.85434, 60.71536, 59.64189, 57.45837, 53.49865,
    50.34034, 49.2573,
  71.53128, 67.44719, 62.60753, 59.70422, 59.70029, 58.85592, 60.74085,
    63.21558, 65.32304, 66.20621, 67.79022, 69.70106, 72.00521, 73.03411,
    72.45726, 72.4124, 72.4092, 72.02244, 71.04708, 70.58475, 69.34588,
    67.23827, 63.83414, 61.61573, 61.20871, 59.88539, 57.93344, 54.25119,
    50.29303, 48.87016,
  71.48013, 68.1069, 64.08553, 60.72916, 60.8099, 58.92272, 59.29606,
    60.57751, 61.64134, 61.93006, 64.13783, 67.30812, 70.84301, 71.81911,
    70.91365, 69.62581, 69.19875, 68.81033, 68.40115, 67.9181, 67.0128,
    65.36415, 63.15838, 61.01101, 60.54426, 59.5718, 58.64468, 56.09729,
    51.6822, 48.84909,
  68.13046, 66.72388, 62.71099, 60.47033, 61.58253, 60.68074, 59.09024,
    58.454, 57.85928, 57.67725, 58.07171, 59.59003, 62.46163, 64.43322,
    63.66306, 62.86469, 61.75833, 61.11706, 61.41788, 62.64576, 62.16327,
    61.01033, 58.86883, 57.1183, 57.09575, 56.51896, 55.60589, 54.50985,
    52.70637, 49.6057,
  53.25108, 54.61431, 55.94336, 56.87229, 58.23757, 59.90253, 58.31375,
    54.97444, 53.80464, 54.06602, 53.73454, 53.23435, 53.06532, 53.68988,
    53.56071, 53.26982, 52.65535, 52.13933, 51.84451, 52.00905, 52.67391,
    53.60006, 53.96588, 53.36357, 53.46157, 53.39155, 52.52992, 50.93831,
    49.75832, 49.19211,
  50.68024, 51.17194, 51.83018, 51.74231, 52.53503, 54.30495, 54.90615,
    52.60572, 50.95472, 51.39385, 51.59251, 51.66992, 51.32209, 51.04238,
    50.85023, 50.38728, 49.69676, 48.78797, 48.69184, 48.72644, 48.58689,
    49.0881, 50.0034, 50.62807, 50.59104, 50.68883, 50.31559, 49.3088,
    48.43719, 47.86386,
  58.45411, 58.71461, 59.00516, 59.34476, 59.60917, 59.85665, 60.06464,
    60.2467, 60.54462, 60.8343, 61.09669, 61.37607, 61.46063, 61.56939,
    61.59621, 61.50764, 61.25467, 60.91069, 60.45352, 59.95393, 59.44809,
    58.9203, 58.63727, 58.58317, 57.09845, 53.56535, 51.24051, 52.96511,
    50.54134, 48.82526,
  58.47339, 58.88183, 59.20447, 59.57188, 59.85907, 60.10663, 60.37376,
    60.6181, 60.90139, 61.14992, 61.37485, 61.58818, 61.70257, 61.69556,
    61.55492, 61.43579, 61.28096, 61.20074, 61.06971, 60.85003, 60.60444,
    60.31079, 60.00001, 59.94705, 59.64028, 58.272, 51.75076, 50.81509,
    50.14135, 49.02345,
  58.42581, 58.84951, 59.25193, 59.64992, 59.88217, 60.18518, 60.49692,
    60.82707, 61.12225, 61.36048, 61.61298, 61.85918, 61.92733, 61.89415,
    61.71025, 61.27356, 60.85363, 60.70834, 60.77262, 60.86946, 61.08523,
    61.22157, 61.187, 61.02459, 60.31122, 59.15102, 58.36694, 53.73978,
    49.42588, 48.93127,
  58.44743, 58.88821, 59.35283, 59.81638, 60.0781, 60.40245, 60.73275,
    61.0167, 61.26002, 61.38706, 61.70486, 62.26722, 62.51572, 62.29162,
    62.16769, 61.90819, 61.3774, 60.77427, 60.54946, 60.7075, 60.98784,
    60.7664, 60.19863, 60.27757, 59.85317, 59.95634, 59.44938, 58.97431,
    58.22894, 50.42899,
  58.47426, 58.88284, 59.37937, 59.79676, 60.08625, 60.56401, 61.09644,
    61.32124, 61.35889, 61.33335, 61.66941, 62.51232, 63.0881, 62.90051,
    62.71624, 62.65537, 62.21385, 61.57602, 61.14497, 60.62717, 60.20567,
    60.00669, 59.69899, 59.9563, 59.80991, 59.44381, 59.52937, 60.45893,
    60.48131, 58.8036,
  58.59267, 58.96845, 59.43118, 59.77116, 60.05926, 60.72079, 61.6831,
    62.24146, 62.24043, 62.20485, 62.43408, 63.10525, 63.71505, 63.34456,
    63.1579, 62.9464, 62.14079, 61.9102, 61.63311, 61.08484, 60.36544,
    59.32819, 59.74218, 59.74475, 59.5763, 59.37365, 59.12366, 59.39261,
    59.45174, 54.1388,
  59.25968, 59.26851, 59.59717, 59.83049, 60.09163, 60.80853, 61.88954,
    62.57064, 62.95742, 63.057, 63.19325, 62.79943, 61.96706, 62.01397,
    61.75174, 61.52692, 61.62514, 60.90123, 59.9968, 59.8167, 59.45342,
    59.32309, 59.52818, 59.78315, 59.73729, 59.59139, 59.71223, 59.66149,
    58.63254, 47.79583,
  61.17883, 60.3599, 60.44448, 60.46865, 60.6134, 61.24215, 61.84384,
    61.07589, 58.68652, 61.23807, 61.49278, 61.69635, 62.00164, 62.25453,
    62.3724, 62.3564, 62.03698, 61.41653, 60.677, 59.91804, 59.37565,
    59.21158, 59.30939, 59.48474, 59.51446, 59.81757, 59.93568, 59.2864,
    58.17902, 47.97482,
  65.17201, 63.63726, 62.58966, 62.08496, 61.8181, 61.63163, 60.76489,
    61.04708, 61.16977, 60.33286, 60.14683, 60.61402, 61.36844, 61.84791,
    62.21901, 62.2691, 62.46843, 62.50467, 62.12849, 61.15695, 60.26009,
    59.62393, 59.2868, 58.91787, 58.98801, 59.7618, 60.01096, 58.81303,
    47.99837, 48.47829,
  69.89088, 69.08509, 67.37684, 65.80633, 64.70822, 63.11005, 61.2111,
    61.59475, 61.58484, 61.45271, 61.12671, 60.56523, 59.58257, 58.98254,
    59.2295, 60.57433, 61.46297, 61.80888, 61.91644, 61.62406, 61.32613,
    60.28912, 59.32549, 58.61162, 58.74937, 59.01316, 58.86754, 53.07859,
    47.93606, 48.03719,
  72.23573, 72.48907, 73.45466, 71.63369, 69.90671, 66.50038, 64.1834,
    62.69997, 62.09554, 62.50493, 61.46355, 60.41239, 60.15248, 57.93094,
    56.19073, 56.50342, 56.58506, 57.39017, 58.98066, 60.65713, 61.10546,
    60.62596, 59.54526, 59.33975, 59.81217, 59.32903, 55.76862, 48.36029,
    48.86276, 48.11701,
  70.70739, 70.37548, 74.02451, 75.76057, 74.76544, 71.19183, 67.46136,
    63.91584, 62.21314, 62.63034, 62.10879, 61.46307, 61.26708, 61.00791,
    60.35476, 59.5013, 59.42758, 58.3822, 57.59951, 58.2058, 60.53709,
    60.49013, 59.39774, 59.23745, 59.52526, 58.76549, 48.6293, 52.70328,
    49.48063, 48.64006,
  62.59777, 64.58605, 66.63924, 69.41885, 71.75043, 71.79614, 66.33279,
    62.23842, 64.42999, 63.22477, 62.90914, 62.40821, 62.51958, 62.43141,
    61.65706, 60.07812, 60.12686, 60.23555, 60.09275, 59.83207, 60.25316,
    60.32952, 59.39849, 57.00472, 56.02628, 57.11291, 48.82742, 50.49826,
    50.25508, 49.2593,
  60.98677, 61.12314, 61.1422, 60.78426, 61.01136, 62.03973, 63.62116,
    64.36916, 62.78272, 63.13464, 63.26634, 62.68774, 62.43433, 62.45356,
    61.73043, 60.73619, 60.34215, 60.6403, 60.79677, 60.05887, 59.77175,
    59.29035, 54.08253, 50.9809, 48.42458, 48.70227, 48.68045, 48.23926,
    48.668, 48.78844,
  61.59479, 61.78101, 61.80736, 61.64079, 61.80869, 62.36299, 63.11331,
    63.27489, 62.83426, 62.44991, 62.137, 61.77981, 61.88722, 61.86303,
    61.58948, 61.48941, 60.75331, 60.64919, 60.47058, 59.39037, 53.6814,
    53.83435, 51.74868, 49.07721, 49.84427, 49.46545, 48.95193, 48.52415,
    48.21626, 48.20781,
  59.06871, 60.73473, 61.29325, 61.3545, 61.58867, 62.34718, 63.08768,
    63.4192, 63.211, 62.7953, 62.6141, 62.48133, 62.48062, 62.7037, 62.02704,
    61.31673, 61.23277, 59.02672, 55.10347, 53.87111, 52.54324, 51.72864,
    49.97422, 49.25933, 49.45699, 49.44051, 48.97311, 48.5294, 48.32182,
    48.26526,
  60.31546, 59.29741, 59.4408, 59.66457, 59.86779, 60.21191, 61.47474,
    62.93391, 63.20068, 63.17049, 63.11712, 63.57153, 64.29914, 64.32013,
    63.5906, 63.346, 63.19944, 61.91992, 58.46328, 55.55479, 52.76686,
    52.2781, 50.74751, 49.70625, 49.85269, 49.68849, 48.87431, 48.25446,
    48.12571, 48.19836,
  66.41998, 63.37588, 60.84857, 60.14064, 60.19247, 59.79596, 59.99412,
    60.8938, 61.85819, 61.84852, 63.13776, 63.58654, 63.86954, 63.91715,
    63.91897, 64.6377, 65.5701, 65.86851, 64.73251, 62.38011, 56.5613,
    53.57197, 51.98853, 51.07535, 50.44428, 49.89797, 49.05202, 48.25106,
    48.10751, 48.13901,
  75.25827, 70.94176, 65.41258, 60.25836, 61.38271, 60.56778, 60.58449,
    60.76251, 60.40124, 60.47694, 60.58828, 59.67177, 58.00491, 57.94751,
    58.4907, 60.65353, 64.33319, 65.9989, 66.09269, 65.11249, 63.09992,
    57.20346, 53.83529, 53.02743, 51.4989, 50.52818, 49.60067, 48.52566,
    48.08865, 48.16598,
  75.60369, 71.98557, 67.21025, 62.58503, 63.41456, 62.95853, 62.83529,
    62.67223, 62.70774, 63.00025, 62.65736, 61.31227, 60.71309, 57.90683,
    55.84964, 55.46582, 56.66457, 59.34445, 61.2947, 61.9491, 61.436,
    58.73544, 55.39079, 54.02399, 52.52205, 51.03223, 50.00221, 48.61544,
    48.06388, 48.16711,
  76.33285, 73.5857, 68.85453, 65.14664, 66.0997, 65.77145, 65.8755,
    65.80175, 65.63309, 65.13737, 63.63785, 62.34103, 62.61458, 61.62761,
    59.80813, 59.09636, 58.80669, 58.84208, 58.71564, 57.43232, 56.99625,
    57.44062, 56.52354, 54.8819, 53.57406, 51.54598, 50.01263, 48.66248,
    48.04136, 48.15074,
  76.07768, 74.35661, 69.73379, 66.80801, 68.52183, 68.44669, 69.00488,
    69.32999, 69.92491, 69.61567, 67.85506, 66.36086, 65.56396, 64.49704,
    63.27758, 62.44261, 61.54638, 60.86659, 59.92504, 58.18887, 56.26261,
    55.72527, 57.27761, 55.54821, 54.70995, 52.48598, 50.44024, 49.03909,
    48.13866, 48.13076,
  75.48134, 74.67163, 69.74332, 66.7205, 69.08225, 69.96018, 70.91833,
    71.73476, 73.25414, 74.02637, 73.82361, 73.75311, 72.93727, 71.90634,
    70.20497, 68.91256, 67.44435, 65.66018, 63.87394, 61.7105, 59.15788,
    57.44369, 57.69876, 56.6121, 56.55614, 54.38415, 51.68602, 49.85959,
    48.78938, 48.25551,
  75.51501, 73.34135, 68.7391, 66.18237, 67.69518, 68.18294, 69.84526,
    72.03391, 74.77351, 76.48687, 77.2459, 78.06565, 78.67357, 78.10365,
    76.59129, 75.46833, 73.80989, 71.99964, 69.49003, 67.20341, 64.95627,
    62.43557, 59.77662, 58.64656, 58.57398, 57.45425, 54.92865, 51.39634,
    49.83355, 48.89075,
  74.98278, 71.90656, 65.20952, 62.10843, 62.75154, 63.06218, 65.57642,
    69.3924, 73.8895, 74.69088, 75.04878, 76.43785, 77.55051, 77.89883,
    76.98248, 76.02004, 74.26475, 72.46972, 70.93391, 68.99317, 66.51084,
    64.1106, 61.24512, 59.42513, 59.47282, 58.44464, 56.64534, 52.9985,
    50.332, 49.37973,
  74.0741, 70.80522, 64.92751, 60.84711, 60.47277, 59.96382, 62.36022,
    66.49727, 69.9352, 70.39033, 71.94571, 74.10465, 75.93256, 76.36497,
    75.40742, 74.66599, 73.34198, 71.38792, 70.24684, 69.30312, 67.39254,
    64.8952, 62.34143, 60.5289, 60.16879, 58.91023, 57.32547, 53.91038,
    50.3482, 49.06595,
  72.03057, 69.12098, 64.0863, 60.44512, 60.37311, 58.85229, 59.61339,
    61.51219, 63.57482, 64.22325, 66.15873, 68.88137, 71.94463, 73.01367,
    71.89336, 70.62556, 69.2285, 67.89089, 67.83304, 67.40452, 65.93398,
    64.02924, 62.27566, 60.63965, 60.10187, 59.20983, 58.19398, 55.68895,
    51.6292, 49.039,
  67.44373, 65.98798, 61.99095, 59.94483, 61.11058, 60.31886, 59.04368,
    58.53606, 58.22447, 58.36702, 59.08057, 60.89762, 63.47823, 65.17233,
    64.8774, 63.76183, 62.33269, 61.39874, 61.8782, 62.7949, 61.86253,
    60.52159, 58.46549, 57.01852, 56.73389, 56.11913, 55.37129, 54.49299,
    52.79364, 49.81316,
  54.61102, 55.51834, 56.46161, 56.99296, 58.46904, 60.03574, 57.97611,
    54.8559, 53.93437, 54.08274, 53.92138, 53.66911, 53.69866, 54.19513,
    54.06861, 53.81174, 53.26221, 52.66658, 52.65882, 52.93306, 53.37451,
    53.94416, 54.09071, 53.52975, 53.5015, 53.07043, 52.37647, 51.00568,
    50.17859, 49.54764,
  51.33446, 51.92634, 52.55931, 52.46385, 53.23616, 54.83834, 55.25356,
    52.93964, 51.48481, 51.94914, 52.10815, 52.2285, 51.80854, 51.45153,
    51.22844, 50.84436, 50.18912, 49.32255, 49.29535, 49.42432, 49.37434,
    49.83764, 50.63207, 51.11912, 51.00813, 51.01957, 50.55546, 49.58865,
    48.91553, 48.40921,
  60.60734, 60.57863, 60.40035, 60.16262, 59.80653, 59.54502, 59.36842,
    59.37664, 59.69257, 60.45154, 61.62553, 62.50701, 62.78076, 63.73011,
    64.5379, 64.91016, 64.96529, 64.86633, 64.52822, 63.9962, 62.79745,
    60.87999, 60.01805, 60.33598, 59.97887, 56.92903, 54.97194, 56.51152,
    53.04073, 51.28395,
  60.4537, 60.13613, 60.17941, 60.12208, 60.00885, 59.96984, 60.06391,
    60.29523, 60.67305, 61.17653, 61.6945, 62.56752, 63.71439, 64.62475,
    65.6929, 67.43747, 69.1028, 71.14375, 73.07249, 74.59402, 75.37347,
    74.83507, 73.6276, 74.38062, 75.01938, 65.31805, 53.21373, 54.84501,
    52.79483, 51.52272,
  60.79137, 60.4874, 60.52021, 60.44096, 60.37922, 60.43546, 60.66238,
    60.98209, 61.3881, 61.82649, 62.35438, 63.09699, 63.39066, 63.50911,
    63.8163, 64.00877, 65.70996, 68.72029, 72.35423, 75.31313, 77.19621,
    78.5872, 79.10796, 79.31844, 78.58484, 73.57497, 64.22865, 55.30761,
    52.02222, 51.6254,
  60.88404, 60.61652, 60.66663, 60.61076, 60.53376, 60.60073, 60.93185,
    61.40243, 62.01038, 62.55176, 63.10426, 63.853, 64.72781, 65.65844,
    66.86905, 66.7832, 65.76485, 66.48967, 69.83469, 74.248, 76.93695,
    78.0126, 76.70779, 79.24836, 77.45401, 75.34947, 75.18392, 67.99656,
    57.72387, 52.45259,
  60.95281, 60.83245, 61.00035, 60.91164, 60.71811, 60.82793, 61.24168,
    61.60543, 62.12872, 62.87769, 63.70584, 64.61461, 65.64618, 66.64074,
    67.80586, 69.34815, 70.66783, 71.53108, 72.8829, 74.79045, 74.17122,
    65.83307, 66.53487, 70.645, 74.21562, 76.67223, 77.36983, 78.09448,
    77.88924, 60.57676,
  60.73148, 60.78077, 61.04434, 61.05222, 60.94206, 61.35406, 62.09887,
    62.36511, 62.33058, 62.48825, 63.19079, 64.52835, 65.99422, 66.81374,
    68.38682, 70.53589, 72.01955, 72.82454, 73.49586, 74.81361, 69.1142,
    62.02748, 65.96815, 67.63227, 70.37345, 74.17668, 78.29073, 78.91709,
    77.75957, 55.00344,
  60.46355, 60.40501, 60.73966, 60.79772, 60.92179, 61.59048, 62.62958,
    63.31275, 63.55956, 63.64632, 63.94834, 64.0441, 64.03758, 64.80991,
    66.08064, 67.37206, 67.69724, 67.21029, 66.6202, 67.0368, 65.24717,
    64.50123, 66.52124, 68.66893, 69.82043, 71.2686, 76.68254, 78.53046,
    70.1973, 50.41049,
  60.71324, 60.2211, 60.49086, 60.583, 60.70502, 61.41679, 62.09627,
    61.52654, 61.55098, 62.22025, 62.82355, 63.61813, 64.62254, 65.03657,
    65.29712, 65.48704, 65.64981, 65.3316, 64.68046, 64.74963, 65.30927,
    66.62959, 68.75122, 70.49969, 70.99581, 74.2271, 78.51176, 77.60788,
    61.52859, 50.60732,
  62.38634, 61.41052, 61.09213, 60.89271, 60.78275, 60.91572, 60.52505,
    61.01409, 61.78381, 62.38183, 63.09043, 63.91698, 64.85583, 66.3648,
    67.9798, 69.11313, 70.12957, 71.10413, 70.98954, 69.3588, 68.36638,
    69.1938, 71.00603, 71.45039, 72.51727, 77.65598, 78.03134, 68.47845,
    50.90138, 51.14072,
  65.49987, 64.59293, 63.62169, 63.04868, 62.81722, 61.96801, 61.06197,
    62.16143, 63.08818, 62.45098, 61.88327, 62.79761, 63.22589, 63.59681,
    64.27686, 66.5271, 68.35571, 69.70519, 70.83497, 72.07865, 73.2963,
    72.32918, 70.49769, 69.50614, 74.70103, 78.05056, 71.34879, 55.47322,
    50.61789, 50.55724,
  69.36806, 68.30487, 69.18109, 67.3614, 66.71872, 65.11275, 64.51796,
    64.40256, 65.30652, 67.20724, 64.23428, 58.94649, 58.06099, 57.72662,
    57.53937, 58.57938, 59.73117, 61.12187, 63.10292, 66.57284, 71.91841,
    73.18404, 71.57686, 74.05656, 77.33929, 73.02345, 57.77878, 50.85248,
    51.3952, 50.60637,
  72.73718, 71.4648, 73.585, 74.07725, 72.07673, 69.45753, 67.46648,
    65.05054, 63.95981, 66.08736, 66.59947, 66.59627, 67.20211, 65.20773,
    62.20041, 59.91865, 60.25214, 60.16508, 60.40092, 62.14224, 66.94319,
    70.05561, 69.9294, 76.00389, 77.66176, 67.76265, 51.31498, 54.69247,
    51.95282, 51.07941,
  65.19491, 66.93646, 68.94218, 70.81825, 72.08199, 70.84686, 65.37951,
    63.28934, 66.12193, 66.56331, 67.42845, 67.55257, 68.71741, 69.22033,
    68.94754, 64.33979, 66.47243, 67.14496, 65.85033, 63.92041, 66.15695,
    68.20844, 66.41135, 61.83757, 61.002, 58.67336, 51.67517, 53.17459,
    52.82309, 51.69096,
  61.16494, 60.94056, 61.29383, 60.78848, 61.07201, 61.97137, 63.88948,
    65.02358, 64.88821, 66.15728, 67.65571, 68.46169, 69.11469, 69.95541,
    69.91087, 69.34949, 69.88123, 72.3314, 74.3428, 72.47652, 68.66005,
    66.30636, 60.00466, 54.2494, 51.25786, 51.62638, 51.2672, 50.97608,
    51.32552, 51.30707,
  63.33519, 63.14068, 62.38187, 61.51414, 61.50679, 62.45865, 63.53352,
    63.89427, 64.44221, 64.63094, 64.84565, 64.88606, 66.88561, 68.25618,
    68.6587, 68.84653, 70.01846, 68.36102, 67.79115, 66.10464, 61.03025,
    58.40132, 53.87721, 52.04387, 52.52338, 52.13966, 51.56635, 51.11892,
    50.79183, 50.74165,
  61.09338, 62.42717, 62.60984, 62.18503, 62.07192, 62.76286, 63.60638,
    64.09016, 64.45132, 64.99072, 64.52295, 63.60033, 63.77034, 65.51494,
    63.71236, 63.10777, 64.16565, 60.81231, 58.42356, 57.12348, 54.82793,
    54.48186, 52.60598, 51.8615, 52.17394, 52.06881, 51.5095, 51.16047,
    50.90937, 50.77164,
  58.52757, 58.37686, 59.19958, 60.24433, 61.49549, 61.85056, 62.66333,
    63.77319, 64.48418, 65.21942, 65.92956, 66.92494, 68.08083, 68.41703,
    66.43208, 64.71082, 62.91679, 61.70184, 59.98946, 57.98484, 54.94961,
    54.74601, 53.13402, 52.19795, 52.36119, 52.29491, 51.35017, 50.79108,
    50.72866, 50.71188,
  62.84283, 60.46622, 58.34053, 58.13445, 58.70024, 59.38088, 60.69164,
    62.61384, 63.40203, 64.06963, 65.39338, 67.15354, 68.54863, 69.63575,
    70.35182, 70.45023, 70.21751, 69.5733, 67.28842, 63.14338, 57.79243,
    55.64365, 54.22192, 53.31433, 52.73476, 52.15984, 51.35479, 50.65766,
    50.63071, 50.64159,
  74.34989, 69.72905, 61.67754, 56.96767, 58.05882, 57.7403, 58.25925,
    59.07443, 59.46925, 60.40384, 61.72683, 61.58778, 60.7384, 61.81528,
    62.96058, 65.44147, 69.76378, 73.83893, 73.91028, 70.98197, 64.86405,
    59.17802, 56.02676, 54.95173, 53.57557, 52.62137, 51.72964, 50.84637,
    50.62937, 50.66558,
  75.33975, 71.02439, 63.70757, 59.01384, 59.54436, 59.22712, 59.51073,
    59.81411, 60.3696, 61.45006, 61.29155, 59.52251, 59.64539, 58.10421,
    57.16473, 57.55379, 59.65568, 63.20416, 65.27821, 65.37782, 64.03143,
    61.03085, 57.69035, 56.01063, 54.57928, 53.07738, 51.99134, 50.99775,
    50.6179, 50.69555,
  77.04834, 73.483, 66.91238, 62.40993, 62.56273, 61.99022, 61.95061,
    61.99165, 62.2104, 62.21397, 60.81008, 59.63606, 60.63089, 60.07921,
    59.03152, 58.90128, 59.44286, 60.49699, 61.20564, 60.52327, 60.3672,
    60.31099, 58.79844, 57.15716, 55.54409, 53.56837, 52.04538, 51.01886,
    50.61788, 50.66418,
  77.65573, 75.31657, 70.02631, 66.81963, 67.50659, 66.73884, 66.68461,
    66.56877, 66.89307, 66.1113, 63.79624, 62.5157, 62.38953, 61.82748,
    61.10806, 60.94247, 60.81009, 61.10566, 61.44027, 61.20834, 60.80614,
    59.76293, 58.77581, 58.12814, 56.77273, 54.41824, 52.48729, 51.41703,
    50.68489, 50.62724,
  77.36595, 75.76501, 70.67699, 68.61277, 69.59691, 69.75735, 70.08007,
    70.56136, 71.60465, 71.95876, 70.38317, 70.51824, 70.06347, 69.03316,
    67.50119, 66.71027, 65.77486, 64.66521, 63.80446, 62.94909, 62.04438,
    60.54043, 58.86272, 58.64542, 58.69563, 56.49935, 53.7857, 52.25765,
    51.26392, 50.70066,
  75.74631, 73.85653, 69.84715, 68.11044, 68.96319, 69.32438, 70.43227,
    72.22935, 74.57011, 75.66936, 76.25076, 77.54721, 78.95537, 79.52163,
    78.46211, 76.86465, 74.78638, 72.19666, 69.80578, 67.62329, 65.64549,
    63.75183, 61.4712, 60.41524, 60.51943, 59.97209, 57.37185, 53.85474,
    52.3623, 51.32993,
  74.2084, 70.85805, 67.01369, 64.92112, 65.22991, 65.36889, 67.92812,
    71.32115, 74.20712, 74.70602, 75.13619, 76.65919, 78.63144, 80.03132,
    79.76153, 78.92265, 76.90322, 74.5612, 72.79627, 70.80765, 68.3952,
    65.96289, 63.12191, 61.41581, 61.53159, 60.91006, 59.37321, 55.57902,
    52.98242, 51.87406,
  72.61579, 69.35593, 65.8134, 63.62558, 62.98603, 62.60959, 65.65442,
    69.79624, 72.3933, 72.938, 74.04705, 75.5932, 77.44197, 78.2507,
    76.98326, 75.97276, 74.99398, 73.20637, 72.29184, 71.50825, 70.04967,
    67.96489, 65.28278, 63.39894, 63.23199, 62.02298, 60.36315, 56.65731,
    52.68433, 51.51692,
  71.68132, 68.78677, 65.757, 62.65713, 62.08929, 60.69878, 62.43715,
    65.43486, 67.37088, 67.7401, 69.43027, 71.65719, 74.0338, 75.01762,
    74.03773, 72.78194, 71.65382, 70.42641, 70.36292, 70.2619, 68.82969,
    67.59563, 66.2278, 64.80334, 64.36283, 63.66051, 62.78761, 59.61699,
    54.21414, 51.31401,
  69.46889, 67.57866, 64.27472, 62.79284, 63.45485, 62.43195, 61.67131,
    61.45094, 61.19231, 61.66994, 62.50718, 64.38995, 66.68725, 67.92189,
    67.73152, 67.27358, 66.0164, 65.355, 65.89381, 66.5247, 65.42294,
    63.56178, 61.47821, 60.47971, 60.48482, 60.2269, 59.67439, 58.89544,
    56.51614, 52.3948,
  57.67789, 58.34168, 58.80876, 59.47752, 61.39578, 63.2997, 61.33264,
    58.02716, 57.02079, 57.50746, 57.30703, 57.08627, 57.01514, 57.29129,
    57.28154, 57.28234, 56.92019, 56.58936, 56.41652, 56.55161, 56.77362,
    57.07774, 56.9315, 56.09828, 56.30193, 56.34209, 55.81268, 54.29254,
    53.3114, 52.33858,
  54.5195, 55.01788, 55.2986, 55.19128, 56.30128, 58.61639, 59.24669,
    56.30173, 54.81898, 55.68171, 56.22838, 56.41378, 55.94061, 55.19772,
    54.62749, 54.13149, 53.31486, 52.26962, 52.26711, 52.36634, 52.20084,
    52.78188, 53.44693, 53.81002, 53.79379, 53.97732, 53.69444, 52.48209,
    51.57917, 50.86472,
  59.21575, 59.54658, 59.90079, 60.44427, 60.87529, 61.54462, 62.14529,
    62.71014, 63.37238, 64.11882, 65.21813, 65.16142, 62.9334, 62.55175,
    62.20271, 61.26408, 60.50818, 60.1736, 59.90687, 60.15874, 59.69163,
    57.77388, 57.72144, 59.10906, 59.86139, 58.12459, 58.43807, 59.8147,
    52.04354, 49.24586,
  63.1539, 63.39159, 62.8546, 63.41898, 63.31416, 63.54142, 64.16409,
    64.85555, 65.65509, 66.66723, 68.1507, 70.01332, 71.29888, 70.43523,
    69.62066, 69.87647, 69.19199, 69.55565, 70.10259, 70.77351, 70.49989,
    69.64371, 68.85315, 70.40223, 70.61958, 64.12931, 55.27865, 57.8484,
    52.13582, 49.94872,
  65.4913, 66.17529, 66.30483, 66.36645, 66.26173, 66.25371, 66.14256,
    66.07451, 66.14597, 66.39358, 66.94983, 68.02347, 69.34679, 71.13712,
    72.20985, 71.19232, 71.9201, 72.57293, 72.19206, 71.91731, 72.09624,
    72.22424, 72.16467, 72.15659, 71.5095, 69.73328, 64.08767, 57.4518,
    51.45935, 50.41355,
  68.44974, 69.50681, 70.66143, 71.71404, 72.31736, 73.03397, 73.07806,
    72.47674, 72.18139, 72.09943, 71.95434, 72.21252, 71.75557, 70.91343,
    72.51231, 73.30472, 71.48004, 71.05366, 72.44422, 72.51772, 72.61176,
    72.3006, 72.38084, 72.91064, 72.34332, 70.86189, 69.39669, 65.19102,
    55.66558, 50.50671,
  71.14404, 71.81001, 73.05991, 73.95633, 74.37806, 74.92532, 75.78303,
    75.83499, 76.3967, 76.18038, 76.13917, 77.07015, 77.53593, 76.90694,
    76.51582, 76.32766, 74.97662, 73.01568, 72.39923, 72.38847, 71.88171,
    70.13692, 71.26756, 72.13676, 72.36442, 71.41579, 70.13924, 70.33922,
    70.17359, 58.91855,
  71.87466, 74.14095, 75.12366, 75.87244, 76.00808, 76.64532, 77.95082,
    78.10052, 77.57161, 77.31006, 77.4598, 78.4089, 79.035, 78.37592,
    78.56676, 78.7014, 77.05984, 74.53317, 72.28941, 71.85802, 71.07333,
    65.44452, 70.05083, 71.68869, 72.02538, 71.58911, 70.99576, 71.4458,
    70.27803, 53.72971,
  70.91414, 74.12546, 75.30118, 76.22962, 76.71395, 77.60965, 79.05139,
    79.45953, 78.93018, 78.53539, 78.20238, 77.46228, 72.32778, 74.1983,
    76.1898, 76.49436, 75.47951, 73.54881, 71.15967, 71.52158, 69.45557,
    68.75517, 71.34113, 72.11491, 72.08718, 71.17587, 71.22768, 71.06709,
    69.26058, 48.33189,
  71.69446, 74.32175, 75.67968, 76.74286, 77.38819, 78.60296, 79.74766,
    79.21603, 76.23003, 77.71831, 76.74229, 75.30685, 74.26737, 74.78114,
    75.07758, 75.76163, 76.14185, 74.86994, 72.02155, 71.11726, 71.34365,
    71.7207, 72.37373, 72.58296, 71.83261, 71.55103, 71.86004, 71.04758,
    63.04914, 48.92333,
  76.18269, 76.81254, 77.1925, 77.64523, 77.68835, 78.12486, 76.6452,
    77.48566, 80.06638, 80.24716, 80.12339, 79.79257, 79.63823, 80.31042,
    80.2579, 78.48809, 78.06453, 77.55352, 76.29381, 74.33442, 72.86005,
    73.00542, 73.83595, 73.32659, 72.06834, 72.62239, 71.69796, 69.8961,
    50.44736, 49.40254,
  79.683, 80.62067, 80.1385, 80.44045, 79.89923, 78.60392, 71.4047, 76.3773,
    75.96645, 77.96987, 79.13006, 78.57889, 77.76506, 77.13, 76.42917,
    77.09515, 77.23932, 76.84964, 76.08915, 75.73058, 75.1966, 73.39529,
    71.82122, 70.45975, 71.01183, 71.73257, 70.31811, 56.50547, 48.83848,
    47.87,
  81.41341, 81.27612, 82.57092, 81.37473, 82.2862, 80.17558, 78.6626,
    78.04493, 78.81826, 79.80041, 75.37156, 64.25363, 62.26188, 62.38559,
    62.50915, 64.31191, 66.02991, 67.25408, 69.04996, 73.38354, 74.79937,
    73.45226, 70.55123, 69.61472, 69.99802, 69.55512, 57.22387, 49.23554,
    49.56943, 48.05497,
  86.09734, 84.37843, 86.38145, 87.28506, 84.99751, 82.58396, 80.3732,
    77.66794, 76.04073, 76.90657, 75.79253, 71.7831, 73.3609, 71.54163,
    64.68174, 64.6862, 64.07034, 64.12714, 64.53983, 67.53975, 73.4717,
    73.20019, 70.48878, 70.73107, 70.48505, 66.54411, 49.76334, 53.41616,
    50.55592, 49.03928,
  83.70898, 85.40009, 87.14161, 88.41821, 88.26501, 86.4, 80.28996, 76.63637,
    78.44093, 77.18156, 77.59773, 77.29356, 77.71827, 77.26347, 74.2209,
    69.94807, 69.79636, 69.83596, 68.64527, 69.48473, 72.32372, 71.80925,
    67.57689, 63.18225, 62.04072, 58.41797, 50.86837, 52.28491, 51.88062,
    49.96517,
  76.19984, 77.40807, 78.02253, 77.25816, 77.16608, 78.22425, 79.84338,
    80.35244, 78.38085, 79.86688, 81.22556, 80.52068, 80.63684, 79.70909,
    77.00858, 74.15966, 72.70032, 72.9007, 73.05466, 72.46412, 71.8467,
    67.70823, 60.93018, 54.67438, 51.33663, 50.96728, 49.77225, 49.2421,
    49.6891, 49.38655,
  76.59315, 76.6934, 77.85168, 77.34803, 77.2316, 78.2245, 81.13638,
    81.94527, 78.99502, 78.35447, 77.31221, 76.27648, 76.17319, 77.04028,
    76.24192, 73.89382, 73.26383, 73.62891, 73.95377, 72.88831, 63.3279,
    60.01859, 54.11208, 52.15548, 52.26055, 51.33002, 50.13102, 49.31616,
    48.66558, 48.40865,
  74.79134, 77.756, 78.62016, 78.76165, 78.91875, 79.92377, 80.75463,
    80.09384, 78.30518, 75.01888, 74.2429, 71.6825, 70.36151, 73.5076,
    71.58287, 70.56378, 71.59347, 68.91488, 67.80833, 63.60228, 56.76924,
    56.4146, 52.67379, 51.50264, 51.74332, 51.29086, 49.82724, 49.3274,
    48.8462, 48.4188,
  67.69566, 68.25661, 70.24359, 72.98869, 75.64079, 77.77444, 79.61707,
    80.92842, 80.61026, 79.15978, 77.42751, 77.49678, 78.41702, 77.1689,
    73.94267, 71.15051, 68.51672, 67.57143, 67.31815, 64.05965, 56.33442,
    56.55655, 53.51717, 51.72209, 51.50745, 51.31823, 49.49423, 48.429,
    48.36205, 48.29687,
  65.94299, 65.81954, 65.34679, 67.20518, 69.37376, 71.87511, 74.60158,
    78.02371, 80.75251, 80.73561, 80.89808, 80.88284, 80.05711, 79.42205,
    77.94701, 77.49406, 77.56165, 77.59057, 75.1525, 68.52625, 58.34351,
    55.97641, 54.0564, 52.84257, 51.19776, 50.31909, 49.55672, 48.1833,
    48.12688, 48.0747,
  76.35802, 71.402, 64.71408, 61.6428, 63.89322, 64.87334, 66.89339,
    69.24806, 70.61093, 73.1349, 76.38712, 75.13477, 71.39603, 73.45226,
    74.55644, 77.55715, 79.86319, 81.51725, 80.4066, 77.43567, 67.9491,
    59.44668, 55.38554, 53.78162, 51.5267, 50.19879, 49.45073, 48.44751,
    48.12225, 48.1053,
  76.50848, 71.61517, 64.96625, 60.91339, 62.31696, 63.03479, 64.34729,
    65.92506, 68.36099, 72.19984, 72.39339, 67.1018, 67.44164, 66.34307,
    65.01846, 64.65108, 67.82542, 73.03321, 76.05584, 75.67827, 70.97389,
    64.11282, 58.01813, 55.14058, 53.17164, 50.96222, 49.70175, 48.60596,
    48.08479, 48.10675,
  77.81966, 73.67094, 66.34754, 62.49755, 62.87661, 63.01835, 63.70827,
    64.81007, 66.8722, 68.71259, 66.20074, 62.87966, 65.6425, 65.50494,
    64.17712, 63.10389, 63.68528, 64.9231, 66.32384, 66.17474, 65.8968,
    65.55579, 62.26384, 58.1343, 54.99483, 51.87402, 49.76427, 48.62511,
    48.04574, 48.11831,
  82.23177, 78.54184, 71.88823, 68.77582, 69.16133, 67.97305, 67.99359,
    68.12018, 70.07793, 70.08693, 65.50887, 63.25399, 64.46236, 64.25882,
    63.36503, 63.02396, 62.57403, 62.51827, 63.1601, 63.89074, 64.35608,
    63.61393, 63.09299, 62.08587, 58.535, 53.22876, 50.21229, 49.14368,
    48.20164, 48.06697,
  85.80301, 84.58763, 77.66445, 75.11973, 77.24063, 77.43103, 76.32948,
    74.74701, 75.72717, 74.44885, 70.45657, 71.03556, 71.25738, 70.67007,
    68.87165, 68.31981, 67.489, 65.00475, 63.42325, 63.15697, 62.9083,
    61.82261, 60.61937, 61.50343, 62.37687, 57.6888, 52.43008, 50.82029,
    49.37293, 48.20726,
  86.31102, 85.18282, 80.59068, 78.80529, 79.52522, 78.88986, 79.92363,
    80.58907, 84.43052, 82.49928, 78.64023, 81.3109, 82.96227, 83.34129,
    80.95918, 79.20067, 77.16975, 73.77039, 69.73254, 67.45242, 65.67543,
    63.85181, 61.9229, 61.38136, 62.74461, 63.03781, 58.85402, 53.57258,
    51.52759, 49.30007,
  86.68903, 83.19039, 76.12872, 73.6037, 73.66399, 73.3297, 75.55608,
    80.45434, 86.1014, 83.17307, 78.93107, 81.53379, 83.45917, 84.34182,
    83.676, 83.06113, 80.86057, 78.37155, 75.99348, 73.45078, 70.47455,
    67.48841, 64.1882, 62.17615, 62.82087, 63.61266, 62.86576, 57.5155,
    53.46917, 50.94051,
  87.72929, 85.41383, 79.62885, 74.7405, 72.78944, 71.7985, 75.64554,
    81.40659, 83.76731, 80.49474, 81.05617, 83.1739, 84.92294, 84.09939,
    81.84213, 81.48985, 80.70433, 79.21443, 78.22984, 76.95422, 75.51972,
    73.37135, 69.52028, 66.61694, 66.53482, 65.46027, 64.28184, 59.31521,
    51.95316, 49.86794,
  85.63642, 82.85806, 78.1539, 74.81582, 73.37097, 70.7149, 73.28813,
    76.23701, 76.4153, 75.42483, 77.56219, 79.79307, 81.43822, 81.14024,
    79.7033, 78.67433, 77.90932, 77.05349, 76.83401, 76.14646, 75.36952,
    75.61921, 74.84165, 72.61639, 72.35811, 71.66785, 71.29383, 67.03757,
    55.44982, 48.9381,
  78.97731, 77.78336, 76.05013, 75.90369, 76.95143, 75.34628, 73.42289,
    71.53282, 68.76852, 69.48027, 70.44073, 72.58708, 74.40613, 74.86073,
    74.50592, 73.63225, 71.90806, 71.06106, 71.97103, 72.59834, 70.266,
    67.30522, 64.83488, 64.16991, 65.12068, 65.58793, 65.82403, 67.06046,
    62.97424, 52.12576,
  66.61009, 67.34935, 67.82333, 68.96024, 73.08679, 76.70291, 72.56055,
    65.20583, 62.78016, 63.55229, 62.98591, 63.08973, 63.57392, 64.02676,
    64.20022, 63.86428, 62.57444, 61.44281, 60.26121, 58.91366, 58.40091,
    58.04145, 56.88389, 55.89777, 56.77742, 57.59643, 57.07968, 55.04219,
    54.56223, 52.521,
  59.42819, 59.99852, 60.06841, 59.50287, 61.74916, 67.10178, 69.01218,
    61.23447, 57.69966, 59.79097, 61.04771, 62.28482, 62.15553, 61.04464,
    59.56512, 58.31525, 55.49204, 52.61019, 52.41393, 52.22194, 51.16787,
    51.72005, 52.27873, 52.46188, 52.9009, 53.78444, 53.66024, 51.63599,
    49.54663, 48.15659,
  50.9379, 51.01993, 51.15727, 51.34136, 51.29688, 51.45785, 51.76698,
    52.18368, 52.72085, 53.60416, 55.63178, 55.60247, 52.08793, 52.25062,
    52.46426, 51.67984, 51.53673, 52.23833, 53.22815, 55.07893, 55.64198,
    53.93597, 54.35166, 56.86549, 58.63248, 58.0141, 62.24174, 64.26168,
    51.50351, 47.59644,
  54.72251, 55.09095, 54.409, 55.23488, 54.61788, 54.26759, 54.71645,
    55.12474, 55.64549, 56.35247, 57.65134, 59.51254, 60.51734, 58.05766,
    56.20185, 56.68007, 55.39008, 56.22978, 57.92635, 59.38895, 58.92812,
    58.02602, 58.28761, 61.79726, 64.64705, 60.79008, 58.43449, 62.56942,
    52.0863, 48.77404,
  53.84082, 54.54028, 55.44203, 56.25694, 56.88462, 57.18473, 57.06408,
    57.19506, 57.51571, 58.01696, 58.65825, 59.77457, 60.9142, 62.49853,
    63.19635, 60.62511, 60.25877, 61.47294, 62.49543, 64.16326, 64.79831,
    65.0183, 65.19208, 65.75751, 65.66488, 64.33259, 64.15932, 61.06427,
    51.60284, 49.69909,
  57.1517, 57.80831, 59.18093, 60.61314, 62.13501, 63.56693, 63.37232,
    62.43882, 62.69367, 63.25554, 63.14796, 63.46488, 62.88554, 61.48917,
    64.37354, 66.00948, 63.14381, 60.42401, 62.81862, 64.87565, 65.33375,
    65.50587, 66.00523, 67.22448, 67.32101, 66.00683, 64.36633, 61.11638,
    53.28598, 48.37201,
  59.47953, 59.24095, 61.34838, 62.89024, 63.95002, 64.15957, 64.17316,
    63.82803, 64.77464, 65.63797, 65.7908, 66.69173, 66.82115, 66.56024,
    66.44524, 66.75552, 66.03003, 63.59591, 64.44151, 64.98115, 65.00233,
    62.71042, 64.57272, 66.46606, 67.50246, 66.33842, 63.92591, 63.92534,
    64.03474, 53.94492,
  61.65852, 63.89696, 67.22997, 68.97461, 68.605, 68.67774, 69.30266,
    68.98154, 68.08056, 67.53885, 67.3972, 67.85061, 68.17889, 67.59016,
    67.93417, 68.82101, 68.22265, 66.11462, 64.29453, 64.63651, 64.45473,
    59.81287, 63.57355, 65.9931, 66.95135, 66.16655, 64.41203, 64.89484,
    64.3494, 51.91499,
  63.35199, 65.59443, 68.38372, 69.04319, 68.45802, 68.40182, 68.63692,
    68.32001, 67.5862, 67.30501, 67.30983, 67.15038, 66.88213, 67.26263,
    67.55801, 67.6913, 67.59232, 66.12984, 64.49968, 64.87772, 63.45119,
    62.94342, 65.42188, 66.73238, 66.83987, 65.21683, 64.80251, 64.71409,
    63.87061, 47.60067,
  63.78024, 66.16979, 69.74118, 69.98277, 69.21026, 69.12724, 69.50958,
    68.54873, 65.49724, 66.93033, 67.24237, 67.09157, 67.43096, 67.98367,
    68.25241, 68.48817, 68.78792, 68.21681, 66.70788, 66.13724, 65.62825,
    65.992, 67.03495, 67.50455, 66.47143, 65.67505, 66.02228, 65.44977,
    61.77352, 47.99283,
  71.80821, 71.99843, 72.06191, 71.56329, 70.21568, 69.92358, 70.06298,
    70.44801, 71.02905, 71.39333, 71.57182, 71.53677, 71.88041, 74.33439,
    75.41222, 72.40021, 72.41357, 72.73133, 72.0414, 69.99947, 68.50649,
    69.44575, 71.00212, 69.99627, 67.55054, 68.26488, 67.0916, 65.17793,
    51.68213, 47.70824,
  77.25786, 78.50759, 77.6573, 77.86508, 75.56573, 73.30112, 71.61772,
    72.08115, 72.07521, 73.338, 74.23177, 74.85006, 74.14629, 72.37514,
    70.62714, 71.80912, 72.38464, 72.17195, 71.64404, 72.66393, 73.31219,
    71.25161, 69.54279, 67.12788, 66.55661, 66.75562, 65.75304, 56.3457,
    47.4617, 45.32185,
  75.0761, 74.53571, 75.88594, 75.01012, 75.14082, 73.31236, 71.71286,
    71.01855, 71.45587, 71.57376, 69.46649, 63.18168, 61.99889, 62.36561,
    63.2307, 65.11298, 66.43419, 66.83009, 67.65491, 68.78366, 70.44334,
    69.61858, 65.28041, 63.58158, 63.78519, 63.63606, 54.01056, 47.96435,
    47.32623, 45.50889,
  80.57586, 78.48132, 81.38655, 81.59654, 78.45669, 75.30724, 72.47144,
    69.23756, 66.66969, 65.67636, 62.62156, 60.58338, 62.88057, 64.31249,
    63.46179, 63.07132, 62.29558, 62.97472, 64.46914, 66.71395, 69.36339,
    68.74613, 64.5505, 64.94914, 64.46384, 59.41942, 48.8021, 50.50064,
    48.82656, 46.69386,
  82.95841, 84.69632, 86.15812, 85.69659, 84.0115, 80.12046, 72.27493,
    68.35732, 68.8653, 66.59657, 66.62238, 65.83581, 66.54836, 67.21262,
    66.62177, 65.70145, 65.90089, 66.16505, 67.187, 69.13435, 68.72688,
    67.36146, 64.50755, 62.8239, 61.506, 55.66136, 49.64001, 50.49632,
    50.50512, 47.79755,
  74.49798, 75.42937, 75.78526, 73.96764, 73.34943, 74.65369, 76.18175,
    75.24993, 71.15096, 70.44476, 70.03662, 67.9016, 68.85182, 69.29456,
    67.4083, 65.94411, 65.69804, 65.94, 66.69998, 67.12, 66.3239, 64.97808,
    61.25669, 55.00671, 51.92659, 50.89275, 48.51733, 47.72336, 48.0911,
    47.08204,
  72.34406, 73.26617, 73.37392, 72.7205, 71.66125, 72.2608, 75.38885,
    74.97952, 71.20436, 69.97025, 68.7748, 67.96173, 68.59277, 68.72506,
    67.78565, 66.92695, 66.34229, 66.94602, 68.19437, 67.87041, 60.46975,
    58.83006, 53.92305, 52.96845, 52.49336, 50.74962, 48.8887, 47.51434,
    46.66593, 46.01974,
  73.15273, 73.68235, 74.1374, 73.57317, 72.35596, 72.25716, 73.78362,
    72.73956, 70.61051, 68.94653, 68.75766, 67.37446, 66.63779, 67.83712,
    66.99145, 66.49098, 66.86711, 67.04706, 67.69187, 66.63757, 55.23716,
    55.61565, 51.99792, 51.18495, 51.5298, 50.80944, 48.61844, 47.72837,
    46.83743, 45.99473,
  69.66998, 67.55288, 68.88592, 70.94205, 71.10037, 70.77667, 71.29453,
    72.38893, 71.62141, 70.33647, 68.22933, 69.04944, 71.12233, 69.24217,
    67.25406, 66.73808, 66.5849, 66.63458, 67.55936, 66.77489, 54.47089,
    56.20054, 53.02122, 51.18865, 50.81407, 50.79139, 48.02192, 46.36592,
    46.22203, 45.8924,
  67.46035, 68.45236, 68.56364, 70.81466, 71.64111, 71.45683, 70.74985,
    70.54597, 70.8337, 69.71549, 70.74635, 72.46137, 71.63348, 69.76596,
    69.67945, 68.31313, 67.14333, 67.30524, 68.51612, 66.95068, 55.89716,
    54.46795, 52.72528, 51.83312, 49.72315, 48.87646, 47.98589, 45.77144,
    45.70479, 45.51725,
  73.86552, 71.41069, 66.78586, 64.69304, 66.92286, 67.23145, 67.71781,
    68.61974, 68.44863, 69.52636, 70.70813, 70.20484, 67.856, 67.66179,
    67.52226, 68.43658, 70.55729, 72.71407, 73.57838, 71.22623, 65.9482,
    57.22022, 53.3632, 51.71511, 49.12804, 47.74014, 47.20711, 46.08861,
    45.66987, 45.52231,
  73.07964, 71.11369, 65.77591, 62.19186, 63.45368, 63.93175, 64.28936,
    65.05883, 67.69128, 70.44188, 70.62595, 67.57466, 66.74518, 65.20927,
    63.92986, 63.87112, 67.34324, 69.27321, 70.2403, 70.09139, 68.22284,
    63.42014, 56.46179, 53.52937, 51.30275, 48.45689, 47.19033, 46.06018,
    45.66922, 45.5382,
  69.50652, 68.10693, 62.81963, 59.97758, 60.41833, 60.78277, 61.13653,
    62.29499, 65.89005, 69.96752, 67.94778, 62.39177, 66.14272, 65.55054,
    63.589, 62.12017, 63.1978, 64.07865, 64.30121, 64.01814, 65.30429,
    66.86838, 62.95317, 58.46691, 54.12249, 49.55318, 47.30915, 46.10518,
    45.65763, 45.54952,
  68.78062, 65.41823, 62.23634, 60.42085, 60.46023, 59.2571, 60.0332,
    60.94565, 65.46413, 67.29987, 60.28568, 56.08381, 58.75273, 59.35056,
    58.9937, 59.50956, 59.37367, 59.64682, 61.23215, 62.05658, 62.00885,
    62.39625, 63.74087, 63.26348, 57.83134, 50.77451, 47.39398, 46.65627,
    45.81538, 45.52087,
  70.46509, 69.61004, 65.47501, 64.26636, 66.6815, 67.6999, 66.70068,
    64.31674, 66.01981, 64.42738, 57.66163, 58.00918, 59.36282, 60.50118,
    59.9815, 61.30484, 61.74288, 59.07819, 58.23808, 58.18449, 57.30874,
    57.04467, 57.13472, 59.72631, 61.94283, 56.11647, 50.27466, 48.7766,
    47.15368, 45.69812,
  76.31982, 75.13859, 72.16587, 73.13283, 72.43999, 69.67542, 71.92524,
    72.74673, 74.43884, 70.24939, 61.96205, 63.75089, 65.47453, 67.34432,
    66.96854, 67.13438, 67.15478, 64.80386, 61.39502, 59.90974, 58.29486,
    57.0732, 56.73777, 57.1092, 59.77943, 62.31186, 58.0465, 51.39099,
    49.32017, 46.70424,
  78.57339, 76.17075, 68.97485, 66.76818, 68.01924, 68.0271, 68.58265,
    71.98531, 76.40669, 74.0368, 65.27798, 66.30111, 66.86178, 67.96397,
    68.58408, 70.27644, 70.23186, 69.43113, 66.83121, 63.56944, 61.34665,
    60.19877, 59.09522, 58.04819, 58.75555, 62.23164, 63.67561, 57.14649,
    52.93024, 49.21367,
  81.09664, 79.48853, 76.03357, 70.90369, 68.63836, 68.09731, 72.59206,
    75.46136, 76.59409, 71.90999, 70.06273, 69.41687, 69.75454, 69.30871,
    68.19884, 70.17034, 72.08141, 72.37409, 71.53362, 69.22972, 67.09521,
    65.96975, 63.11029, 60.36602, 60.72532, 61.85601, 64.02072, 59.30364,
    51.27424, 48.26603,
  80.98975, 78.91241, 75.47762, 71.24522, 69.94242, 67.26675, 71.8654,
    74.39576, 70.90638, 69.28156, 70.69458, 70.15937, 69.60106, 69.67673,
    70.75034, 72.16081, 73.33721, 73.13802, 72.77354, 72.05127, 71.12498,
    70.97514, 70.53973, 69.41659, 68.68134, 68.24413, 68.23466, 66.60377,
    54.70826, 46.20265,
  79.47055, 76.16611, 75.76386, 74.59163, 75.47243, 75.00159, 74.32706,
    71.6466, 66.01993, 67.76791, 68.42966, 68.33477, 68.27075, 68.71655,
    70.46651, 71.18715, 70.65833, 71.40021, 71.53439, 71.67278, 70.55596,
    69.37914, 68.67565, 68.37132, 68.40462, 67.97852, 67.44626, 67.64838,
    66.17651, 50.61524,
  70.41817, 71.22266, 72.53221, 72.43471, 73.9558, 75.24968, 74.27679,
    68.52621, 64.57116, 65.56889, 65.16885, 65.89964, 66.53481, 66.40946,
    66.98842, 66.82875, 65.26963, 63.95387, 61.89596, 58.20424, 56.03444,
    55.15536, 53.22551, 52.34373, 54.30335, 56.57119, 57.30383, 55.85307,
    55.77332, 51.68024,
  66.86559, 67.60515, 67.80348, 67.54057, 70.49558, 72.77256, 73.05428,
    69.87477, 63.06828, 65.94606, 68.07294, 68.87663, 68.27269, 66.97414,
    64.9733, 62.60495, 58.03961, 53.63297, 52.98668, 51.80491, 49.73119,
    49.78326, 49.84502, 49.91399, 50.72525, 52.38517, 52.99318, 50.75352,
    47.83951, 45.55374,
  45.23001, 46.01266, 46.63243, 47.3441, 47.92778, 48.55965, 49.16097,
    49.80699, 50.48327, 51.14795, 52.534, 52.51272, 50.33348, 50.19815,
    49.4574, 47.79467, 46.78643, 46.57569, 46.80172, 47.96715, 48.45229,
    47.39941, 47.71175, 48.62257, 48.73513, 47.62457, 49.74772, 49.49328,
    40.57339, 37.87613,
  53.72097, 54.72719, 54.86104, 56.05467, 56.40386, 56.81841, 57.64846,
    58.46648, 59.2468, 59.84747, 60.4919, 61.44446, 61.75692, 59.51557,
    57.24954, 55.66763, 53.08575, 52.32866, 52.53112, 52.81261, 52.21907,
    51.21362, 51.08683, 53.52106, 56.64714, 54.21332, 50.70538, 51.32437,
    41.69794, 38.86592,
  56.51199, 57.69432, 58.61637, 59.75887, 60.82781, 61.9774, 63.1761,
    64.46353, 65.25765, 65.3148, 65.36025, 65.5583, 65.66843, 65.79929,
    65.71208, 64.19247, 62.38418, 61.76252, 61.17734, 61.32687, 62.446,
    63.36094, 62.86478, 62.72113, 63.51321, 61.11385, 56.46119, 50.66502,
    42.26097, 40.03352,
  61.92437, 63.55574, 65.06134, 65.71374, 65.96513, 66.33408, 66.61406,
    66.69109, 66.83302, 66.72285, 66.49579, 66.80794, 66.88498, 66.39202,
    66.5794, 66.62731, 65.76604, 64.26707, 64.17699, 64.76823, 65.29261,
    65.21686, 62.80838, 65.97495, 66.30006, 63.90824, 58.99171, 49.72215,
    42.44083, 38.6195,
  65.97199, 66.01431, 66.22079, 66.41119, 66.35939, 66.60309, 67.12725,
    67.29597, 67.37212, 67.17382, 66.95294, 67.28017, 67.40923, 67.16558,
    66.86987, 66.69959, 65.94834, 64.4936, 63.81278, 65.27359, 65.49883,
    62.18554, 62.07028, 64.65169, 65.97618, 64.98641, 59.28039, 59.12578,
    54.46577, 42.0671,
  66.86403, 67.08007, 67.314, 67.43482, 66.91707, 66.98779, 67.71951,
    67.74376, 67.35694, 67.10954, 67.06161, 67.5217, 67.83669, 67.17362,
    66.79686, 67.51527, 68.17107, 66.62563, 65.00472, 64.99592, 63.60989,
    59.29438, 60.13626, 61.55986, 64.09969, 62.48269, 60.01388, 63.05054,
    62.01984, 40.37897,
  67.45712, 67.59975, 67.71688, 67.66239, 67.19419, 67.23503, 67.68333,
    67.61124, 67.03827, 66.72225, 66.5416, 66.22092, 65.79116, 65.62106,
    65.71705, 66.44621, 66.72554, 65.61378, 61.98296, 61.45726, 59.20021,
    57.74925, 58.47374, 60.98609, 61.01896, 57.68885, 59.76343, 63.21549,
    55.28086, 37.87383,
  67.83264, 67.91971, 68.02512, 68.0823, 67.56595, 67.50806, 67.87083,
    67.40374, 66.86503, 66.80167, 66.74483, 66.63637, 66.4395, 66.37281,
    66.52504, 66.70615, 66.6917, 65.97259, 61.36066, 60.33725, 59.02969,
    58.88453, 60.91785, 62.16903, 58.99157, 57.43178, 62.55836, 60.21972,
    46.94387, 38.21051,
  70.85441, 70.98798, 71.02177, 70.88156, 70.27069, 70.35049, 70.46945,
    70.80687, 71.29723, 71.28727, 71.18674, 71.05408, 70.99498, 72.03301,
    72.28231, 70.19676, 69.78793, 69.89877, 69.37638, 68.0133, 67.10471,
    67.60149, 68.44393, 67.50913, 64.08666, 63.48997, 62.29452, 53.68389,
    41.25992, 37.87312,
  77.30634, 77.7543, 77.73638, 78.1312, 76.62585, 74.5308, 73.68369,
    74.22417, 74.29065, 74.6599, 74.88804, 75.31662, 74.83464, 73.21748,
    71.51063, 71.41553, 70.96767, 70.09187, 68.74814, 68.07012, 67.89133,
    66.957, 64.58032, 59.96645, 63.14295, 65.3855, 59.51319, 42.198,
    38.01067, 36.47531,
  77.17981, 77.46096, 78.83415, 78.58958, 79.90842, 78.29321, 76.47868,
    75.48287, 74.84988, 75.05473, 74.62293, 69.99489, 69.35808, 68.72391,
    68.2233, 67.80452, 67.4983, 66.80701, 64.09177, 61.34259, 62.46061,
    58.5952, 51.11995, 47.58072, 48.75046, 47.88151, 41.915, 37.77254,
    37.36549, 36.46364,
  78.56063, 75.22551, 77.64913, 79.12901, 78.42331, 76.8709, 75.5301,
    72.41882, 69.32191, 69.07726, 68.23212, 67.07467, 67.23714, 67.62376,
    66.73521, 65.8351, 61.87998, 58.84325, 56.46469, 55.76629, 56.81161,
    53.03714, 46.53857, 51.55051, 53.88718, 42.75008, 37.8187, 38.38442,
    37.84694, 36.94504,
  84.70306, 84.98124, 85.8968, 86.49562, 85.28336, 81.75857, 74.29489,
    70.65157, 71.44972, 68.99554, 69.67848, 69.07653, 69.02579, 69.01236,
    67.75095, 66.27097, 64.82944, 61.21614, 58.50193, 59.35223, 57.57761,
    50.7643, 47.31336, 48.18734, 48.53305, 41.34302, 38.5806, 38.71392,
    38.70349, 37.46732,
  76.40472, 76.88971, 77.01733, 75.43235, 74.41383, 74.15737, 74.34506,
    74.79135, 72.19893, 71.92401, 72.46526, 70.72687, 71.84032, 72.24454,
    69.92668, 67.73835, 66.4866, 66.11176, 66.03522, 65.65229, 56.69152,
    50.72894, 50.41081, 43.6195, 40.30636, 39.51621, 38.13033, 37.58946,
    37.75898, 37.223,
  70.61259, 70.82553, 70.73928, 70.46476, 70.44828, 71.65217, 75.24635,
    76.27854, 73.41846, 72.98997, 72.37173, 71.62397, 71.47587, 70.74881,
    69.42752, 67.39283, 66.30772, 66.02695, 66.48167, 64.08786, 51.15251,
    48.27816, 42.89388, 40.77815, 39.63663, 39.06244, 38.03881, 37.38934,
    37.05786, 36.71546,
  73.03072, 73.52209, 73.77605, 73.57731, 73.45156, 74.3202, 75.08511,
    74.5288, 73.63131, 72.57243, 71.99982, 70.34963, 69.42716, 69.57678,
    67.98394, 66.78954, 66.1931, 61.6791, 58.57493, 54.44188, 44.40686,
    43.46108, 41.23458, 40.33192, 39.61297, 38.84961, 38.02279, 37.51732,
    37.09206, 36.6776,
  72.22783, 72.16972, 72.19006, 72.30489, 72.83686, 72.76463, 73.26825,
    73.86171, 73.18302, 72.33401, 70.95132, 70.93249, 71.67801, 69.61019,
    67.7232, 66.54449, 63.15256, 57.41719, 57.53577, 55.09946, 43.16376,
    43.28387, 41.51811, 40.24632, 39.25685, 38.94154, 37.90714, 37.02858,
    36.87961, 36.6709,
  70.13849, 70.64697, 70.52905, 70.80947, 70.82875, 71.1397, 71.34039,
    71.72219, 72.05971, 70.99983, 70.9971, 71.29003, 70.31628, 69.25665,
    68.39573, 66.37325, 58.5588, 53.76236, 55.96667, 52.65641, 43.63885,
    42.6202, 40.98669, 39.84026, 38.39708, 38.05201, 37.61166, 36.72673,
    36.6197, 36.4962,
  72.22428, 71.23137, 69.77388, 68.94243, 69.35651, 69.28232, 69.73767,
    70.35972, 70.18019, 70.04607, 70.53334, 69.89101, 68.54294, 68.79589,
    68.41862, 68.19434, 68.7785, 69.28771, 69.4761, 63.66444, 51.74745,
    44.45892, 40.86638, 39.80971, 38.01084, 37.48245, 37.25693, 36.78484,
    36.60199, 36.48886,
  71.83494, 70.67893, 69.28696, 68.40289, 68.85284, 69.17291, 69.66831,
    70.00661, 70.19704, 70.78908, 70.66294, 69.24672, 69.02787, 68.73243,
    68.19942, 67.73017, 66.35641, 65.80725, 64.94119, 62.96368, 56.0587,
    48.02374, 42.20472, 40.51165, 38.87491, 37.80181, 37.25385, 36.83842,
    36.59369, 36.48346,
  71.2162, 70.25758, 68.59994, 67.65813, 67.97923, 68.28868, 68.58297,
    68.77264, 69.01513, 69.28847, 68.54106, 67.46175, 67.53327, 67.24668,
    63.76376, 58.98501, 56.50494, 55.56322, 56.0574, 55.19188, 53.33117,
    51.31157, 46.48228, 42.52259, 39.98356, 38.39201, 37.30993, 36.86928,
    36.5888, 36.48317,
  71.66824, 69.85547, 68.25774, 67.13247, 67.24854, 67.13941, 67.21869,
    67.20234, 67.59383, 67.51228, 64.51364, 62.17689, 62.45535, 60.44471,
    57.15746, 54.02077, 51.47801, 50.21323, 49.85232, 49.294, 50.10702,
    50.71593, 49.27032, 48.10807, 43.68335, 39.42011, 37.43405, 37.09538,
    36.63641, 36.47797,
  71.67315, 70.08929, 68.31255, 67.17639, 67.45057, 67.40331, 66.94432,
    65.64435, 65.4901, 63.40942, 59.37475, 59.52072, 59.53195, 58.2187,
    55.38495, 53.11819, 51.06656, 48.32829, 47.03762, 46.61543, 47.31419,
    47.92923, 46.09316, 46.53304, 46.18158, 41.80575, 38.28071, 37.91938,
    37.18069, 36.5546,
  73.91934, 72.61603, 71.27062, 70.35671, 70.1503, 69.7504, 69.80453,
    69.99365, 70.2793, 67.34309, 63.16444, 64.56074, 64.6958, 63.43594,
    60.24662, 56.86134, 54.1464, 51.12599, 48.14576, 47.2178, 47.54119,
    47.06887, 45.38269, 44.4475, 44.6046, 44.50674, 41.3791, 38.72552,
    37.96959, 36.92889,
  75.86434, 76.28911, 73.48731, 72.23273, 72.11903, 71.77442, 71.65968,
    72.16465, 73.06904, 71.96719, 66.99339, 68.01215, 67.39275, 64.95516,
    61.44225, 58.11457, 54.54974, 52.10785, 49.34495, 47.10581, 47.19848,
    46.85495, 45.18478, 43.7689, 42.74291, 43.80354, 43.97407, 41.20198,
    39.57914, 37.97716,
  78.35784, 79.1311, 76.83599, 74.97557, 74.07822, 73.35313, 73.74992,
    74.52726, 74.27317, 71.87424, 69.83724, 69.75949, 68.58301, 64.55013,
    59.6548, 56.4292, 53.96534, 52.04827, 50.04421, 48.0674, 48.17723,
    47.89228, 45.37768, 43.43684, 42.92063, 43.139, 44.08392, 42.4879,
    39.22491, 37.73468,
  78.62272, 79.01708, 76.63631, 75.01619, 74.54233, 73.75663, 74.02104,
    74.24524, 73.57118, 71.00224, 70.72692, 70.46364, 68.75851, 64.99516,
    60.92923, 57.51094, 55.17002, 53.9366, 52.60001, 51.43578, 52.90959,
    54.71116, 53.29811, 49.75279, 47.35434, 46.72889, 47.41251, 46.15265,
    40.04067, 36.72192,
  78.39046, 78.5505, 76.89172, 76.10527, 76.35178, 75.8536, 75.23134,
    74.57409, 73.6003, 73.39333, 73.14944, 73.10777, 72.19613, 69.03796,
    65.8805, 62.46074, 59.4649, 58.14486, 57.5105, 57.11134, 57.45984,
    56.24891, 52.75259, 50.18953, 48.55633, 47.92806, 47.25226, 48.55102,
    45.61353, 38.48083,
  73.98461, 74.17814, 74.91423, 75.3707, 75.7135, 75.98436, 75.01031,
    73.08101, 72.27797, 72.12859, 71.60458, 71.08594, 70.6199, 70.26141,
    68.32648, 64.83631, 61.73421, 59.52909, 56.23475, 52.56004, 51.06801,
    49.30056, 47.11703, 45.47354, 45.08871, 44.89514, 44.12171, 42.52161,
    41.93219, 39.41615,
  71.2754, 71.40401, 71.6566, 71.67553, 72.25346, 73.3914, 73.31525,
    71.32209, 70.06705, 70.19887, 70.1215, 69.77088, 69.03043, 68.11183,
    65.22414, 59.80874, 54.41053, 49.9922, 47.97067, 45.87429, 44.07509,
    43.30925, 42.62835, 41.94801, 41.60235, 41.68558, 41.24659, 39.72849,
    38.03444, 36.6782,
  38.00857, 38.0952, 38.1963, 38.35655, 38.42174, 38.51331, 38.62879,
    38.81765, 39.02848, 39.23848, 40.17945, 40.313, 38.97288, 39.23704,
    39.47263, 39.22093, 39.27851, 39.56013, 39.87642, 40.74376, 41.30789,
    40.74794, 40.87804, 41.73891, 42.29671, 41.84882, 43.98195, 45.13567,
    39.94281, 38.31733,
  40.26813, 40.45903, 40.22422, 40.6464, 40.54489, 40.44491, 40.66005,
    40.8644, 41.08655, 41.3392, 41.69636, 42.34795, 42.89571, 42.1528,
    41.77015, 42.13527, 41.7414, 42.11876, 42.82839, 43.45943, 43.54494,
    43.3092, 43.5226, 44.66196, 48.68797, 49.35691, 43.86637, 45.96446,
    40.49565, 38.87411,
  41.99858, 42.12512, 42.22738, 42.40677, 42.53799, 42.68571, 42.8205,
    43.01579, 43.27638, 43.53421, 43.83111, 44.4155, 44.91485, 45.7034,
    46.18612, 45.4693, 45.6263, 46.28679, 46.62134, 47.17664, 48.49162,
    50.08851, 50.59356, 49.68991, 52.86371, 54.53905, 46.87103, 45.35263,
    40.56803, 39.55027,
  45.54598, 45.847, 46.28656, 46.76184, 47.18579, 47.76767, 47.87529,
    47.64535, 47.87006, 48.23713, 48.33819, 48.69904, 48.7077, 48.24187,
    49.51948, 50.67896, 49.73368, 48.40775, 48.89661, 49.59797, 51.6944,
    52.15862, 50.15524, 54.53793, 56.34484, 50.01566, 49.18415, 44.49569,
    40.76675, 38.77466,
  49.32145, 49.14281, 49.56858, 50.05282, 50.27064, 50.22609, 50.2703,
    50.26377, 50.8051, 51.21808, 50.88625, 50.93642, 51.00341, 51.25124,
    51.53666, 51.96551, 51.132, 49.38796, 49.3351, 54.15041, 55.89894,
    47.89523, 48.16173, 49.57499, 51.53335, 50.86006, 47.35819, 47.74631,
    47.06211, 40.91568,
  52.16354, 52.7917, 53.85316, 55.12582, 54.89797, 54.39596, 54.96116,
    55.21575, 55.01374, 55.37606, 55.94141, 57.92817, 60.19591, 59.60458,
    58.95599, 67.31365, 76.14036, 61.63567, 52.20518, 52.72541, 50.16349,
    46.919, 47.67242, 48.9031, 51.13105, 50.05833, 53.27656, 67.82219,
    59.24355, 39.51443,
  56.61951, 57.84317, 59.15714, 60.42083, 60.44699, 60.37645, 61.42183,
    62.71635, 62.02829, 60.78154, 59.96637, 57.7286, 54.9139, 54.77893,
    58.44431, 63.32818, 59.38172, 52.82245, 49.70467, 49.25635, 47.78721,
    46.81697, 47.38936, 49.63999, 50.46326, 47.24072, 54.65688, 68.14849,
    54.75875, 37.95312,
  58.75283, 59.64875, 60.53704, 61.1552, 60.04705, 60.54634, 61.19434,
    56.85161, 53.62001, 52.84385, 51.52526, 50.06551, 48.9604, 49.13471,
    49.83673, 50.56322, 50.88027, 50.10318, 47.61458, 47.0753, 46.29493,
    46.14186, 47.68408, 49.47123, 48.40693, 46.47975, 55.16668, 58.78534,
    43.65789, 38.60468,
  60.13731, 60.05363, 60.24868, 59.47358, 58.0334, 57.8399, 55.10314,
    53.52212, 53.89808, 53.81986, 53.2317, 52.61824, 52.43105, 56.17884,
    58.65914, 53.61664, 52.87801, 54.35648, 54.12642, 50.97601, 48.70116,
    50.89706, 55.01019, 54.68444, 49.65047, 49.89757, 52.07967, 48.70881,
    40.50071, 38.39141,
  67.8401, 67.65842, 67.61557, 67.59109, 66.88554, 63.62594, 57.80481,
    58.98254, 59.16031, 60.62703, 62.27362, 64.98373, 65.04298, 62.1684,
    58.70882, 59.62701, 60.04819, 59.19863, 56.74206, 55.10783, 55.33593,
    54.62817, 53.51839, 49.82372, 56.64848, 69.30046, 56.5125, 41.02328,
    38.57398, 37.47963,
  72.49349, 71.61314, 71.31815, 70.23947, 69.76219, 69.23284, 68.43158,
    68.33473, 68.63511, 70.11413, 71.39933, 61.4355, 57.76417, 57.19149,
    56.82936, 56.78149, 56.89791, 55.81142, 53.99227, 52.72651, 54.1607,
    52.26021, 47.26652, 44.22129, 45.78011, 46.83368, 42.01238, 38.32251,
    38.01569, 37.41741,
  79.12325, 74.6218, 77.45826, 77.72676, 76.53533, 74.39521, 72.68095,
    69.18667, 66.10782, 66.53274, 64.32567, 58.12542, 59.33389, 58.73923,
    54.49423, 54.15771, 52.18633, 50.87943, 49.33971, 48.82463, 50.23894,
    48.34864, 43.07057, 47.89527, 50.75752, 40.8754, 38.14383, 38.54941,
    38.33966, 37.73247,
  85.6746, 85.13545, 86.60751, 85.64673, 83.5061, 78.53603, 70.14952,
    66.2594, 66.78217, 65.00646, 65.49034, 63.62389, 64.39938, 64.50597,
    56.83229, 52.66935, 50.98275, 49.74508, 48.31426, 49.53496, 49.75238,
    46.0631, 43.12501, 46.28321, 47.91914, 39.98986, 38.59069, 38.72509,
    38.80735, 38.05998,
  78.39889, 79.87823, 78.45849, 75.53738, 73.11365, 72.18522, 72.59471,
    71.93899, 68.92611, 67.85719, 68.52032, 67.49432, 69.74155, 73.23728,
    76.52563, 63.00985, 52.99868, 54.05732, 54.18567, 53.25001, 48.66161,
    47.73281, 50.35605, 42.97709, 40.10101, 39.37255, 38.51549, 38.14242,
    38.31353, 37.9357,
  69.30502, 68.7213, 68.08052, 67.19734, 66.66293, 68.79956, 74.09669,
    73.38357, 69.63618, 68.71618, 67.69505, 67.18752, 67.93864, 71.28321,
    72.41407, 58.34627, 56.50175, 54.09328, 54.83625, 55.87987, 51.93416,
    46.31165, 41.45043, 39.85888, 39.28391, 39.24117, 38.52489, 38.03819,
    37.81461, 37.59472,
  67.43951, 67.19063, 67.30325, 66.89768, 66.61697, 67.22033, 67.91117,
    67.45668, 66.52927, 65.65344, 65.81359, 62.5828, 59.16735, 60.00832,
    57.02909, 54.60196, 53.3241, 50.052, 49.33215, 47.97869, 42.40139,
    41.22422, 39.68626, 39.24546, 39.2841, 39.09156, 38.56982, 38.12716,
    37.82179, 37.56213,
  66.83799, 66.24351, 65.9566, 65.68076, 65.75946, 65.28047, 65.42865,
    66.0149, 65.26589, 63.49651, 59.12776, 58.8079, 61.22271, 57.01949,
    53.69485, 51.57643, 49.50937, 47.12755, 48.18741, 47.24868, 40.64659,
    40.98944, 40.08489, 39.24547, 38.99564, 39.13571, 38.50092, 37.83393,
    37.70013, 37.56421,
  64.38889, 63.42784, 61.85334, 61.33655, 60.63522, 60.55583, 60.18433,
    59.96048, 59.7552, 57.18173, 57.58302, 59.28363, 57.2936, 55.98452,
    55.86595, 51.68948, 46.99421, 44.68465, 46.92731, 45.97822, 40.96396,
    40.87971, 40.14989, 39.44765, 38.66624, 38.58744, 38.28104, 37.65279,
    37.56609, 37.47355,
  62.42216, 60.35358, 57.42773, 55.69549, 55.33257, 54.5806, 54.2767,
    54.24164, 53.31789, 52.7386, 54.41008, 53.43601, 49.45299, 50.26609,
    50.72799, 50.30056, 50.91861, 51.74183, 53.75465, 52.44313, 46.52342,
    42.38915, 40.13057, 39.61002, 38.50198, 38.1606, 38.02097, 37.67695,
    37.5369, 37.46085,
  58.88385, 56.81592, 54.21612, 52.0281, 51.55696, 51.16613, 50.9597,
    50.83346, 50.94862, 53.02696, 53.44981, 49.73456, 49.32643, 49.8464,
    49.84131, 49.39919, 50.25592, 51.37708, 52.02768, 52.02482, 48.84115,
    44.20012, 40.70029, 39.94376, 38.98323, 38.29121, 37.99365, 37.7218,
    37.53265, 37.45902,
  56.42146, 54.74336, 52.37892, 50.53054, 49.92551, 49.74882, 49.72285,
    49.82454, 50.61102, 52.37383, 50.99663, 48.24543, 49.47524, 49.71007,
    48.79163, 47.37903, 46.83759, 46.44383, 46.69113, 46.31727, 45.44455,
    44.79839, 42.84983, 40.98463, 39.57164, 38.6511, 38.01448, 37.71882,
    37.53361, 37.45873,
  56.73292, 54.08742, 52.08805, 50.69344, 50.14458, 49.3155, 49.24186,
    49.06057, 50.33822, 50.86852, 47.96807, 46.21068, 46.76868, 46.50294,
    45.69743, 44.93659, 44.07507, 43.47123, 43.29115, 42.83268, 44.35852,
    45.42348, 43.45641, 43.79549, 41.64723, 39.29238, 38.05907, 37.8386,
    37.57243, 37.45547,
  55.75907, 54.20304, 51.94302, 50.56918, 50.83456, 50.73119, 49.80712,
    48.26123, 48.19017, 47.11289, 44.30256, 44.00629, 44.33965, 44.45382,
    44.01236, 44.14003, 44.02314, 42.70896, 42.06437, 41.73296, 42.7063,
    43.36485, 41.39611, 42.55433, 42.89287, 40.53364, 38.53449, 38.36037,
    37.90919, 37.50502,
  55.82686, 54.50797, 53.35826, 52.57324, 51.95454, 50.94728, 50.71339,
    50.04764, 49.97677, 47.10123, 43.90372, 44.63653, 45.30168, 45.88691,
    45.72913, 45.40523, 45.19337, 44.08885, 42.44155, 41.66974, 41.65037,
    41.55086, 41.04161, 40.95846, 41.58043, 41.93043, 40.30662, 38.77941,
    38.35783, 37.72142,
  55.23234, 55.35086, 52.5854, 51.36696, 51.27144, 50.57619, 49.53036,
    49.18342, 50.21835, 48.06563, 44.62379, 45.50233, 46.25417, 46.51002,
    46.33382, 46.17767, 45.39642, 44.73336, 43.4607, 41.96974, 41.88195,
    41.97167, 41.53119, 40.78412, 40.29624, 41.3253, 41.62494, 40.0899,
    39.26727, 38.3126,
  57.01915, 58.20304, 56.55233, 53.96762, 52.17235, 51.02124, 51.52916,
    52.05661, 50.23907, 47.46319, 46.13081, 46.76222, 47.4363, 46.77048,
    45.66029, 45.36752, 44.99759, 44.56263, 43.71686, 42.44012, 42.4558,
    42.56849, 41.39713, 40.47226, 40.45734, 40.81879, 41.75057, 40.9888,
    39.10616, 38.11225,
  58.50279, 58.73205, 55.52162, 53.38088, 52.39216, 51.00042, 51.60774,
    51.30959, 48.38382, 46.39225, 46.37737, 46.79974, 46.88587, 46.21962,
    45.52866, 45.00329, 44.54892, 44.36372, 43.85572, 42.97034, 43.58127,
    45.00904, 45.06186, 43.66426, 42.7543, 42.67838, 43.74767, 43.39867,
    39.62796, 37.51209,
  57.87461, 56.96453, 54.76554, 53.89869, 53.67162, 52.38148, 51.54106,
    49.58096, 46.36254, 45.95158, 45.86275, 46.24846, 46.56624, 46.37894,
    46.50547, 46.23751, 45.63742, 45.64038, 45.8962, 46.03709, 46.54081,
    46.45452, 45.15033, 44.04322, 43.39768, 43.40675, 43.42608, 44.76867,
    43.07498, 38.5972,
  55.43422, 54.01986, 54.18718, 54.55828, 54.47866, 54.67986, 52.46078,
    48.09238, 45.96721, 46.0046, 45.55236, 45.71833, 46.34708, 47.23061,
    48.29287, 48.73794, 48.63559, 48.55229, 47.32262, 45.51637, 44.93563,
    44.11163, 42.91224, 42.06891, 42.0111, 42.16027, 41.93416, 41.14886,
    41.01282, 39.24897,
  55.3036, 54.9569, 54.47625, 53.51665, 53.47939, 55.36401, 55.59534,
    50.93952, 47.98539, 48.8778, 49.65077, 50.44592, 50.71484, 50.75925,
    50.39703, 49.417, 47.48698, 45.36634, 44.30309, 43.03355, 41.9436,
    41.46307, 40.99512, 40.56201, 40.36484, 40.50509, 40.24051, 39.37103,
    38.51137, 37.63908,
  34.41295, 34.45992, 34.51171, 34.56678, 34.57142, 34.59274, 34.64426,
    34.71805, 34.82654, 34.96165, 35.73571, 35.85794, 34.81732, 34.93778,
    35.06995, 34.80795, 34.76669, 34.88663, 35.01793, 35.67567, 36.04379,
    35.49647, 35.48247, 36.14775, 36.61637, 36.32289, 38.37555, 39.51841,
    36.06237, 34.93421,
  35.30495, 35.39688, 35.16482, 35.43977, 35.34047, 35.21943, 35.3275,
    35.44881, 35.5504, 35.69313, 35.97344, 36.46432, 36.82853, 36.16573,
    35.83158, 36.00666, 35.61444, 35.83006, 36.38461, 36.91142, 37.00872,
    36.69418, 36.87481, 37.69219, 41.65337, 42.59907, 38.38747, 40.46236,
    36.67566, 35.39382,
  35.87669, 35.95721, 35.96561, 36.04602, 36.06992, 36.11911, 36.18385,
    36.27992, 36.40704, 36.48421, 36.57258, 36.91302, 37.20658, 37.73478,
    37.98868, 37.36044, 37.44008, 37.9493, 38.24394, 38.71748, 39.82655,
    41.14459, 41.76965, 41.07739, 45.22084, 47.59921, 40.57039, 40.13347,
    36.71649, 35.8946,
  37.47121, 37.68396, 37.96407, 38.26969, 38.57305, 39.0771, 39.24352,
    39.06413, 39.16301, 39.31143, 39.23093, 39.48244, 39.39651, 38.9583,
    39.98281, 40.99894, 40.39912, 39.59021, 40.09268, 40.74463, 42.7493,
    43.49805, 41.79591, 46.20676, 48.20926, 42.81705, 42.52087, 39.37217,
    36.68876, 35.3444,
  40.17329, 40.15577, 40.53837, 40.9551, 41.12746, 41.24334, 41.42946,
    41.42319, 41.77071, 41.84558, 41.33924, 41.20778, 41.17865, 41.37608,
    41.79689, 42.30402, 41.66151, 40.81273, 40.92509, 45.55437, 47.07527,
    40.53329, 40.54131, 41.75531, 43.40587, 42.68927, 40.36366, 40.65325,
    40.88777, 36.84246,
  42.25892, 42.78672, 43.56451, 44.51997, 44.25375, 43.79604, 44.30501,
    44.48119, 44.18813, 44.23703, 44.29585, 45.68606, 47.3363, 47.11777,
    46.1889, 54.39051, 63.051, 50.94879, 43.24837, 44.24025, 42.35892,
    39.46544, 39.90624, 40.66993, 42.77397, 41.85047, 45.92464, 60.06942,
    52.61498, 35.8403,
  44.85564, 45.81577, 46.86648, 47.97301, 48.20382, 48.39674, 49.70423,
    51.17566, 50.97647, 50.34552, 49.98544, 48.34725, 46.25429, 45.8315,
    50.199, 56.18916, 51.9076, 44.5592, 42.04165, 41.62452, 40.38116,
    39.60855, 40.02481, 41.85378, 42.9062, 40.13078, 49.64577, 64.55004,
    49.92892, 34.68319,
  48.10984, 49.2522, 50.4253, 51.55849, 51.38233, 52.53857, 53.8743,
    51.15377, 48.6314, 47.76327, 46.39836, 44.52821, 42.91958, 42.43927,
    43.0267, 43.62214, 43.13463, 42.24004, 40.53946, 40.1755, 39.60726,
    39.41536, 40.59451, 42.17606, 41.68066, 39.72804, 50.05122, 54.44281,
    39.57975, 35.58508,
  51.8222, 52.23577, 52.74335, 52.45917, 51.67521, 51.74524, 49.6232,
    47.91019, 47.47153, 46.64082, 45.41169, 44.01896, 43.03307, 45.59917,
    47.15257, 43.40234, 43.00831, 44.20036, 44.16368, 41.95615, 40.3063,
    41.89521, 45.44091, 45.46061, 41.96897, 41.99525, 46.83773, 45.95818,
    37.40507, 35.37831,
  56.20378, 57.67955, 57.50978, 57.52762, 55.88889, 51.51624, 47.02502,
    47.3665, 47.12358, 47.26024, 48.05872, 50.38058, 50.64042, 48.72459,
    46.19378, 46.49698, 47.00161, 46.69529, 45.47183, 45.34174, 45.86712,
    46.17848, 46.1053, 43.65032, 50.29175, 60.7979, 50.77605, 38.2199,
    35.65569, 34.45675,
  80.83257, 80.23926, 74.46548, 64.10169, 61.97561, 58.50232, 54.51573,
    55.80727, 56.54286, 65.04108, 70.66231, 50.02303, 45.58144, 44.90227,
    44.71247, 45.73228, 46.51001, 46.19566, 44.94037, 44.62173, 47.04002,
    46.30397, 42.23582, 39.51398, 42.10283, 44.26504, 39.22218, 35.20195,
    34.91573, 34.36473,
  85.52544, 81.88111, 85.39519, 86.30402, 85.97726, 75.73618, 72.9323,
    64.68514, 54.37793, 56.91019, 55.15254, 45.52738, 47.19905, 47.88556,
    45.00322, 45.32893, 44.12999, 43.46058, 42.40197, 42.46468, 45.07085,
    43.57531, 38.58989, 42.84459, 44.8442, 37.23665, 34.86913, 35.30352,
    35.19789, 34.61356,
  91.0792, 92.18233, 96.11959, 96.44221, 95.63686, 91.88626, 81.27127,
    57.14009, 58.56019, 54.34, 53.22348, 47.82845, 50.94222, 52.75495,
    46.78902, 44.75971, 43.86695, 42.70191, 41.49073, 43.28309, 44.39499,
    41.14776, 38.36433, 42.5262, 43.79269, 36.58121, 35.21051, 35.43678,
    35.68716, 34.91839,
  90.01815, 94.71539, 93.49185, 90.58638, 87.69466, 84.7413, 82.17343,
    82.54183, 81.70971, 77.67587, 82.72838, 77.84803, 76.9995, 74.09904,
    65.3012, 52.14144, 44.11625, 45.67833, 46.69556, 47.05577, 43.43553,
    42.84066, 44.78258, 39.343, 37.0279, 36.01177, 35.22448, 34.92559,
    35.25237, 34.83669,
  76.50202, 75.68814, 71.74802, 68.9158, 66.64011, 79.04524, 84.57434,
    85.2785, 82.35302, 81.92549, 79.97086, 63.06026, 53.60103, 60.6001,
    62.17834, 48.44401, 47.95125, 47.03582, 50.07821, 51.24227, 45.8594,
    41.93583, 38.36883, 36.44609, 35.88494, 36.04176, 35.30549, 34.84832,
    34.74294, 34.52755,
  62.48341, 61.28895, 60.97417, 60.50585, 61.06841, 64.72889, 68.04577,
    65.48835, 62.12918, 58.29402, 55.27124, 51.15009, 47.58174, 50.1194,
    48.63625, 46.95861, 47.15682, 44.93498, 45.73185, 44.91817, 39.08444,
    37.45609, 35.97142, 35.71506, 35.96362, 35.90994, 35.42728, 34.93582,
    34.7062, 34.48079,
  58.89295, 57.6357, 56.87175, 56.51887, 56.61301, 55.90841, 55.26111,
    54.73997, 53.89212, 53.17501, 49.00116, 48.83935, 52.09138, 48.85701,
    46.20802, 45.36678, 44.21933, 42.33933, 44.63337, 43.63196, 36.68513,
    37.1343, 36.5185, 35.74424, 35.63623, 35.92184, 35.3642, 34.70379,
    34.59526, 34.46058,
  54.65888, 54.30035, 53.12862, 52.6194, 51.99568, 52.06218, 51.65575,
    51.43087, 51.19553, 48.59055, 48.54627, 50.60964, 49.29162, 48.4017,
    49.43403, 46.41095, 42.05629, 39.94913, 43.36529, 42.49066, 37.14872,
    37.32612, 36.79857, 36.05233, 35.32834, 35.48191, 35.12972, 34.524,
    34.45617, 34.37746,
  53.74393, 52.66161, 50.45203, 49.1264, 48.89556, 48.2998, 48.05137,
    48.04047, 46.97207, 45.91436, 47.64959, 46.62997, 42.28395, 42.82676,
    43.43174, 43.023, 43.68236, 44.70855, 47.79493, 46.77814, 41.06514,
    38.30991, 37.02224, 36.3325, 35.28628, 35.06544, 34.89825, 34.534,
    34.4188, 34.36143,
  51.84005, 51.20711, 48.85415, 46.91321, 46.54068, 46.13103, 45.76693,
    45.30425, 44.80759, 46.49438, 46.47844, 42.13199, 40.61309, 40.8207,
    40.80193, 40.48906, 42.026, 44.06443, 45.86353, 46.72078, 44.0162,
    40.17219, 37.52264, 36.65319, 35.74422, 35.15342, 34.86195, 34.5705,
    34.40637, 34.35544,
  49.93108, 49.10328, 47.06624, 45.31937, 44.71986, 44.42848, 44.0878,
    43.70186, 44.00299, 45.50351, 43.38814, 39.94236, 40.74738, 41.14479,
    40.64383, 39.82817, 39.91244, 40.20848, 41.29992, 41.66768, 41.26085,
    40.87637, 39.4534, 37.58855, 36.18201, 35.40337, 34.86112, 34.56932,
    34.42338, 34.37236,
  49.37367, 47.40342, 45.7153, 44.60685, 44.06768, 43.4186, 43.36597,
    43.12829, 44.47277, 44.85465, 41.46786, 39.47675, 40.13833, 40.03807,
    39.48972, 39.01735, 38.44009, 38.20536, 38.34229, 38.19294, 39.78444,
    40.69196, 40.16325, 40.67379, 38.4613, 36.03596, 34.9458, 34.70311,
    34.47207, 34.37943,
  48.10162, 47.01592, 45.07996, 44.11086, 44.81969, 45.36597, 45.07874,
    44.08528, 44.51119, 43.17659, 39.65736, 38.84976, 38.94648, 38.90756,
    38.45987, 38.69878, 38.69402, 37.67617, 37.29472, 37.19236, 38.39481,
    38.84638, 37.74271, 39.31818, 39.76857, 37.24731, 35.31491, 35.19492,
    34.78614, 34.43081,
  48.25286, 47.27627, 46.55503, 46.36565, 46.38728, 46.33101, 46.66307,
    46.47088, 46.77226, 43.29922, 39.15686, 39.11609, 39.37202, 39.80969,
    39.73404, 39.7059, 39.87285, 39.04573, 37.70033, 37.24491, 37.48331,
    37.45077, 37.07225, 37.28329, 38.36321, 38.7389, 37.07577, 35.62055,
    35.19207, 34.60638,
  48.56265, 49.16692, 46.71493, 45.95352, 46.24748, 46.01574, 45.35649,
    45.34829, 46.63806, 43.51976, 39.12059, 39.39272, 39.96446, 40.1991,
    40.30273, 40.415, 40.07016, 39.8715, 38.66911, 37.2775, 37.51847,
    37.78065, 37.51926, 36.83083, 36.37928, 37.66972, 37.9859, 36.56286,
    36.0388, 35.07999,
  49.62758, 51.28588, 49.99189, 47.90523, 46.30737, 45.31655, 46.2678,
    47.36136, 45.71568, 42.24252, 40.0353, 40.33545, 41.11544, 40.59692,
    39.73035, 39.73616, 39.70711, 39.75047, 38.99458, 37.71297, 38.14652,
    38.46915, 37.23021, 36.3601, 36.34333, 36.83972, 38.14465, 37.43699,
    35.89197, 34.90936,
  50.42477, 51.3483, 48.48751, 46.78635, 45.95939, 44.96407, 46.31116,
    46.71186, 43.67995, 41.10569, 40.43095, 40.62821, 40.80577, 40.23716,
    39.69339, 39.35986, 39.14667, 39.2876, 38.78819, 37.75168, 38.70621,
    40.57531, 40.67434, 39.05727, 38.19868, 38.3156, 39.83718, 39.67392,
    36.23228, 34.36987,
  49.72509, 49.40635, 47.64819, 47.20586, 47.53747, 46.9398, 46.99329,
    45.32524, 41.82842, 40.76055, 40.0951, 40.18024, 40.32669, 40.09854,
    40.2423, 39.92815, 39.28446, 39.40126, 39.70988, 39.72992, 40.99994,
    41.5679, 40.44065, 39.12385, 38.52828, 38.75049, 39.02834, 40.90135,
    39.4094, 35.33657,
  47.39241, 46.3489, 46.84928, 47.8735, 48.74672, 49.85167, 48.09315,
    43.85659, 41.38604, 40.68796, 39.3717, 38.76993, 38.84377, 39.59364,
    40.84767, 41.34621, 41.45018, 41.90759, 40.85552, 39.32737, 39.20973,
    38.70221, 37.70378, 37.11305, 37.2518, 37.70263, 37.77875, 37.40564,
    37.84855, 35.9673,
  46.75497, 46.70509, 46.58953, 46.07419, 46.48332, 49.15805, 49.82726,
    45.00412, 41.72645, 41.74281, 41.77597, 42.08494, 42.2891, 42.86782,
    43.22588, 42.83815, 41.50917, 39.97241, 39.0288, 37.81399, 36.99955,
    36.70362, 36.424, 36.24741, 36.27785, 36.66487, 36.6223, 35.98972,
    35.37296, 34.57327,
  27.18716, 27.22879, 27.26296, 27.29217, 27.29062, 27.29332, 27.32204,
    27.38622, 27.46734, 27.58602, 28.57875, 28.65001, 27.52222, 27.7324,
    27.84934, 27.49991, 27.41833, 27.4807, 27.55809, 28.2473, 28.60331,
    27.99621, 27.92228, 28.5323, 28.90293, 28.52145, 30.99784, 32.56301,
    29.20949, 27.93506,
  27.76056, 27.80093, 27.55374, 27.83155, 27.68151, 27.54731, 27.62172,
    27.69508, 27.78328, 27.96567, 28.32717, 28.91177, 29.32718, 28.59758,
    28.24017, 28.31861, 27.81604, 27.92375, 28.49895, 29.10174, 29.06034,
    28.52411, 28.56021, 29.44736, 33.30561, 33.71862, 31.1887, 34.08117,
    30.05143, 28.58759,
  27.82901, 27.86639, 27.82856, 27.88075, 27.87264, 27.85616, 27.8948,
    27.96904, 28.03543, 28.07676, 28.19915, 28.62971, 28.96764, 29.57927,
    29.78399, 28.93853, 28.88113, 29.33983, 29.48936, 29.86248, 30.96249,
    32.33658, 32.98437, 32.47831, 36.70699, 38.74545, 33.51337, 33.6268,
    29.93744, 29.07658,
  28.50375, 28.56274, 28.77843, 28.97958, 29.256, 29.79464, 29.89902,
    29.58492, 29.5806, 29.7759, 29.80082, 30.14605, 30.00685, 29.61624,
    30.71708, 31.84991, 31.15955, 30.1336, 30.49096, 31.0566, 33.53277,
    34.56055, 33.14833, 37.51849, 39.03126, 35.2237, 35.81717, 32.99484,
    29.90334, 28.34013,
  30.31503, 30.08878, 30.3743, 30.75195, 31.03158, 31.21028, 31.22793,
    31.00446, 31.33384, 31.45633, 31.02546, 30.92401, 30.85542, 31.19387,
    31.8811, 32.47255, 31.8154, 30.95949, 31.3319, 36.09012, 37.2742,
    31.7394, 31.63529, 33.20646, 35.13722, 34.74404, 32.93493, 33.79488,
    34.66413, 30.10407,
  31.9522, 32.23416, 32.9687, 33.93417, 33.80293, 33.39298, 33.61822,
    33.30429, 32.51702, 32.19962, 32.06262, 33.72219, 35.8154, 35.86438,
    35.47456, 43.34237, 50.64926, 40.6926, 34.10824, 35.71014, 33.68796,
    30.37617, 30.85284, 31.80704, 34.48191, 33.90145, 37.42915, 50.16181,
    44.47142, 29.31833,
  34.03738, 34.65054, 35.52605, 36.59404, 36.79639, 36.73482, 37.82542,
    39.06121, 38.45451, 37.68028, 37.62116, 36.60458, 35.19982, 35.40576,
    40.339, 46.70124, 43.43081, 35.85835, 33.1666, 32.89437, 31.47423,
    30.48483, 31.07537, 33.54053, 34.96685, 32.60447, 42.52185, 56.34388,
    42.87714, 27.8952,
  36.4183, 37.32895, 38.60258, 39.93225, 39.92342, 41.81396, 43.8643,
    40.92916, 38.02779, 37.0229, 35.85617, 34.21233, 32.89619, 32.81818,
    34.2362, 35.2917, 34.52598, 33.35757, 31.6144, 31.30259, 30.71853,
    30.5046, 31.99528, 34.41207, 34.02474, 32.50718, 44.59057, 48.69827,
    33.47635, 28.27132,
  40.33382, 41.10454, 42.29804, 42.59201, 42.57444, 43.57552, 41.67484,
    39.28014, 38.18806, 36.87453, 35.21212, 33.5547, 32.54737, 35.92824,
    37.95762, 34.13689, 33.76657, 35.3096, 35.46561, 32.96754, 30.99012,
    32.84799, 37.59734, 38.19201, 34.28723, 34.87616, 40.35696, 38.2289,
    30.25621, 28.18953,
  45.1833, 47.38105, 48.78318, 50.23124, 49.14212, 44.07942, 38.88898,
    38.18501, 36.78771, 35.55074, 35.91482, 38.88511, 40.14152, 38.85797,
    36.66305, 36.83465, 37.50644, 37.91098, 36.34302, 34.84262, 35.23352,
    36.03665, 36.89069, 34.95305, 41.3091, 51.53924, 42.57724, 31.02816,
    28.5831, 27.39781,
  62.09985, 64.34018, 58.40017, 51.20633, 49.254, 47.36509, 42.91496,
    43.75215, 44.66486, 52.17664, 55.27932, 39.08245, 35.17446, 34.77916,
    34.31987, 34.97992, 35.95713, 35.97192, 34.86774, 34.76336, 37.28027,
    36.76413, 33.59483, 31.4554, 35.06506, 38.18181, 32.62857, 28.19117,
    27.83636, 27.26769,
  76.81833, 64.55352, 69.31398, 71.07466, 68.15092, 58.16465, 58.27846,
    52.5167, 44.18169, 47.38983, 45.59695, 33.90945, 35.34697, 36.35888,
    34.36755, 34.70766, 33.89842, 33.63785, 33.21244, 33.69248, 36.5994,
    35.25705, 30.91005, 35.03545, 36.79031, 30.05175, 27.74371, 28.17406,
    28.11074, 27.50227,
  90.67171, 91.71152, 96.49803, 97.91159, 98.94431, 91.9247, 68.15115,
    47.06377, 45.67271, 42.42172, 39.97241, 34.04671, 38.21724, 40.29668,
    35.83625, 34.67931, 34.29402, 33.50051, 32.69183, 34.80118, 36.22011,
    33.28241, 30.58586, 35.57136, 36.64267, 29.3842, 28.02091, 28.30945,
    28.61939, 27.77932,
  93.82462, 100.061, 99.88773, 97.8175, 87.07053, 76.54108, 73.89113,
    70.00063, 60.67797, 57.06768, 63.76006, 59.88167, 60.16986, 58.61168,
    51.7122, 41.65384, 34.7179, 36.25348, 37.57025, 38.4905, 35.41172,
    34.79731, 36.44482, 32.34538, 30.0818, 28.76064, 28.04744, 27.81867,
    28.22389, 27.70334,
  68.88299, 71.93655, 65.95624, 60.91376, 55.44648, 64.33645, 88.09031,
    86.31239, 77.06507, 76.0272, 70.14292, 53.77902, 43.69955, 48.82643,
    50.80676, 38.50586, 38.49363, 38.36159, 42.01007, 42.89001, 38.03658,
    34.70704, 31.41235, 29.19408, 28.53277, 28.7957, 28.11932, 27.69736,
    27.67944, 27.42961,
  52.821, 50.72538, 49.51402, 48.50959, 49.33854, 54.77656, 60.66777,
    58.7489, 54.76784, 51.17445, 47.1571, 40.26114, 36.54558, 39.84058,
    39.71539, 37.94593, 38.92538, 37.22917, 38.71396, 37.92215, 32.31455,
    30.29099, 28.65517, 28.49217, 28.78458, 28.67056, 28.23769, 27.80764,
    27.61952, 27.35654,
  48.41356, 46.86258, 46.35725, 46.65569, 47.77269, 48.07388, 47.71843,
    46.89827, 44.71888, 42.16422, 37.91133, 37.79471, 41.80061, 39.62128,
    37.5686, 37.33877, 36.55429, 34.91307, 37.06891, 35.56685, 29.27835,
    29.6818, 29.2895, 28.6426, 28.53174, 28.70211, 28.17576, 27.57597,
    27.50491, 27.34677,
  45.29065, 45.43346, 45.04699, 45.33232, 45.08925, 45.00764, 44.18325,
    43.07144, 41.69567, 38.26885, 37.91937, 40.64802, 40.32547, 39.89946,
    41.23402, 38.7305, 34.53815, 32.4113, 35.76118, 34.51385, 29.70115,
    30.08503, 29.7645, 28.98996, 28.18104, 28.33002, 27.96036, 27.40245,
    27.35136, 27.26687,
  46.40702, 46.23966, 44.33368, 43.11262, 42.7616, 41.9754, 41.16461,
    40.18829, 38.13903, 36.24018, 38.19332, 38.0329, 34.08456, 34.92543,
    35.7638, 35.15876, 35.55946, 36.50724, 39.47043, 38.22984, 33.16152,
    31.03917, 30.00139, 29.19149, 28.12101, 27.93355, 27.77785, 27.41226,
    27.32095, 27.24489,
  46.10609, 45.38789, 43.24979, 41.35372, 40.93966, 40.38716, 39.53172,
    38.19316, 36.68186, 37.66504, 37.72221, 33.71913, 31.94628, 32.31,
    32.24044, 31.87336, 33.61757, 35.99715, 38.08978, 38.72468, 36.23012,
    32.82374, 30.34738, 29.45051, 28.55656, 27.99308, 27.72942, 27.43699,
    27.31006, 27.24776,
  44.40562, 43.84149, 41.92479, 40.31199, 39.79014, 39.39169, 38.48041,
    37.04894, 36.22805, 37.0304, 34.54704, 30.96337, 31.67123, 32.18438,
    31.82179, 31.269, 31.6373, 32.31849, 33.69416, 34.23445, 34.02761,
    33.61117, 32.09996, 30.22069, 28.96914, 28.25063, 27.72207, 27.43047,
    27.32508, 27.24968,
  44.11127, 42.64508, 41.06835, 39.97729, 39.38916, 38.50517, 37.61122,
    36.20509, 36.36234, 35.86396, 32.12132, 30.28844, 31.27514, 31.49918,
    31.19102, 30.93326, 30.57769, 30.54696, 30.7891, 30.76671, 32.09942,
    32.71187, 32.70251, 33.02219, 31.08656, 28.81886, 27.81732, 27.56652,
    27.37627, 27.26329,
  42.96688, 42.0962, 40.24051, 39.22381, 39.60961, 39.69246, 38.66974,
    36.74208, 36.34048, 34.24387, 30.59607, 30.15015, 30.67236, 30.80464,
    30.48266, 30.8881, 30.85296, 29.96135, 29.65885, 29.64411, 30.75644,
    30.99628, 30.44086, 32.03613, 32.43247, 29.8764, 28.15242, 28.04668,
    27.64887, 27.30261,
  42.20784, 41.5847, 40.87136, 40.59731, 40.608, 40.46069, 40.26027, 39.2909,
    38.65766, 34.42392, 30.36292, 30.67384, 31.26761, 31.80362, 31.74673,
    31.85736, 32.0725, 31.16692, 29.96582, 29.74172, 30.00583, 29.94467,
    29.69955, 30.02484, 31.30324, 31.48475, 29.7017, 28.40713, 28.04331,
    27.44303,
  41.98885, 42.62402, 40.71972, 40.30322, 40.71001, 40.42726, 39.43831,
    38.71106, 38.83959, 34.62856, 30.3856, 30.9591, 31.8068, 32.21891,
    32.44531, 32.63493, 32.34557, 32.0168, 30.77729, 29.61942, 29.92988,
    30.17689, 29.96942, 29.28206, 29.0567, 30.36375, 30.4772, 29.14027,
    28.85873, 27.84715,
  42.69133, 44.81192, 44.20403, 42.41998, 40.89246, 39.71809, 40.12982,
    40.17692, 37.52187, 33.33433, 31.06861, 31.74657, 32.76406, 32.46717,
    31.88006, 32.00861, 31.92797, 31.94772, 31.11891, 29.93171, 30.46416,
    30.6946, 29.5423, 28.76725, 28.78706, 29.38246, 30.67234, 29.8689,
    28.7121, 27.67765,
  44.08259, 45.73437, 43.14617, 41.44767, 40.60165, 39.44512, 40.10476,
    39.4435, 35.27145, 32.03074, 31.45505, 32.14393, 32.62877, 32.17327,
    31.71577, 31.4806, 31.29794, 31.49298, 30.92628, 29.88662, 30.88921,
    32.52716, 32.44033, 31.01988, 30.44051, 30.64992, 32.31277, 31.99321,
    28.86446, 27.19122,
  43.60479, 43.79181, 41.98196, 41.60371, 42.11198, 41.4383, 40.97347,
    37.98127, 33.29364, 31.64647, 31.24529, 31.81365, 32.20494, 31.9725,
    32.13216, 31.86182, 31.20903, 31.30571, 31.50988, 31.54168, 32.99726,
    33.44906, 32.3751, 31.09594, 30.77839, 30.99998, 31.44857, 33.41758,
    31.68025, 27.97547,
  41.21791, 40.50715, 41.0009, 42.21153, 43.62709, 44.7713, 42.24105,
    36.71058, 32.99937, 31.69376, 30.52725, 30.26229, 30.47656, 31.16919,
    32.31681, 32.82812, 32.92273, 33.4384, 32.38651, 31.08685, 31.19028,
    30.75313, 29.79949, 29.27696, 29.5346, 30.08693, 30.24503, 30.13876,
    30.72101, 28.56754,
  40.17265, 40.33743, 40.43192, 40.30531, 41.08055, 43.8325, 43.53608,
    37.24799, 32.92383, 32.39143, 32.46895, 32.87276, 33.25208, 33.94534,
    34.33891, 34.18145, 33.04905, 31.82114, 30.92058, 29.73838, 29.0998,
    28.89612, 28.69369, 28.61832, 28.72262, 29.28279, 29.30722, 28.73249,
    28.26845, 27.4502,
  23.86898, 23.8971, 23.93814, 23.95028, 23.9353, 23.9499, 23.9574, 23.96959,
    24.04285, 24.10741, 24.98634, 24.96228, 24.09548, 24.28953, 24.38354,
    24.09521, 24.01023, 24.0285, 24.04863, 24.6015, 24.82294, 24.2864,
    24.19791, 24.71475, 25.02395, 24.6349, 26.90487, 28.09933, 25.50202,
    24.45684,
  24.27038, 24.24596, 24.0521, 24.28745, 24.16296, 24.03496, 24.06882,
    24.12893, 24.20557, 24.35204, 24.70778, 25.25916, 25.5912, 24.88036,
    24.63233, 24.608, 24.1838, 24.24378, 24.64379, 25.08, 25.02318, 24.48705,
    24.49465, 25.14324, 28.71606, 28.75038, 27.44785, 30.20073, 26.53227,
    25.0566,
  24.18623, 24.18607, 24.14021, 24.19198, 24.16513, 24.12547, 24.1251,
    24.20562, 24.29365, 24.32489, 24.45022, 24.87734, 25.14263, 25.61879,
    25.65392, 24.87295, 24.77479, 25.0993, 25.18674, 25.36104, 26.11077,
    27.20572, 28.00246, 27.42964, 31.76377, 33.66748, 29.82344, 30.01608,
    26.61166, 25.6223,
  24.24987, 24.26151, 24.45457, 24.61137, 24.83909, 25.28658, 25.31948,
    25.08337, 25.15408, 25.35324, 25.37353, 25.76483, 25.60125, 25.25733,
    26.12651, 27.02145, 26.27483, 25.43208, 25.68827, 26.03419, 28.25031,
    29.2266, 28.23337, 32.27988, 33.40524, 31.2602, 32.37805, 29.60238,
    26.57946, 24.98216,
  24.84026, 24.65126, 24.88366, 25.23753, 25.50665, 25.65771, 25.70154,
    25.56131, 26.04861, 26.27406, 26.05503, 26.03458, 25.95389, 26.18647,
    26.7812, 27.32247, 26.51762, 25.88834, 26.25482, 30.72146, 31.53806,
    27.26854, 27.22647, 28.88101, 30.4607, 30.34528, 29.48131, 30.40435,
    31.08108, 26.48739,
  25.18218, 25.33045, 26.05599, 26.98012, 26.75949, 26.32225, 26.5729,
    26.3681, 25.96779, 26.0123, 25.99651, 27.81783, 29.72438, 29.87043,
    29.242, 36.62861, 42.42663, 33.99295, 28.95894, 30.83532, 29.04864,
    26.10124, 26.5894, 27.26718, 29.99457, 29.54323, 32.8408, 43.77356,
    38.88543, 25.91232,
  25.87023, 26.24816, 27.02953, 27.88674, 27.86284, 27.58907, 28.67886,
    30.07909, 30.08319, 30.06195, 30.55514, 30.07774, 29.29975, 29.47843,
    34.28267, 40.60691, 37.8779, 30.73847, 28.47629, 28.22743, 26.95995,
    26.10718, 26.73125, 29.14168, 30.48362, 28.3298, 37.71333, 49.77474,
    37.78806, 24.60662,
  26.86563, 27.35781, 28.38777, 29.40701, 29.31446, 31.26465, 33.41637,
    31.35679, 29.65734, 29.59818, 29.41441, 28.42933, 27.63067, 27.67464,
    29.54522, 30.73007, 29.61666, 28.26824, 26.98962, 26.80743, 26.35877,
    26.18158, 27.56879, 29.93667, 29.53089, 28.16198, 40.03418, 43.13841,
    29.93303, 24.78234,
  29.40467, 29.90511, 31.07836, 31.32602, 31.80033, 33.19926, 31.96186,
    30.25004, 29.915, 29.59701, 28.82913, 27.91202, 27.29596, 30.43233,
    31.75993, 28.6083, 28.69453, 30.12335, 30.19713, 28.02776, 26.40277,
    27.99786, 32.3267, 32.64918, 29.42531, 29.93399, 36.11372, 33.98682,
    26.79415, 24.75911,
  33.10424, 34.88399, 36.42192, 37.57895, 37.61973, 33.79853, 29.71511,
    29.30623, 28.77633, 28.10974, 29.06977, 31.98848, 33.59838, 33.09718,
    31.47798, 31.54246, 32.25471, 32.74564, 31.32941, 30.05686, 30.17706,
    31.12811, 32.23335, 30.69958, 36.30072, 44.68606, 37.41823, 27.66176,
    25.2317, 24.11652,
  45.0151, 47.5119, 43.85041, 38.8681, 37.95148, 36.07644, 32.30973,
    33.49494, 34.71312, 42.14206, 44.50444, 32.74622, 30.1017, 29.70902,
    29.11338, 29.99102, 31.08467, 31.10932, 30.04962, 30.12661, 32.60275,
    32.48681, 29.45553, 27.55419, 31.59645, 35.1403, 29.40215, 24.90015,
    24.47545, 23.99033,
  57.71826, 47.64993, 50.41352, 52.41971, 50.16653, 43.946, 45.32436,
    41.12631, 35.0323, 39.29753, 38.38062, 28.24906, 29.46583, 30.27259,
    29.02083, 29.33904, 28.88368, 28.82407, 28.4196, 29.12847, 32.33902,
    31.16512, 27.16827, 30.7938, 32.02616, 26.54717, 24.48074, 24.79421,
    24.71913, 24.15806,
  66.46813, 65.2419, 82.75854, 86.41251, 83.88375, 73.02731, 55.05316,
    37.93839, 35.9649, 34.35471, 32.05408, 27.28113, 31.66502, 33.94335,
    30.39145, 29.62252, 29.60417, 28.82042, 28.23021, 30.48858, 32.18106,
    29.55957, 26.85873, 32.10592, 32.65664, 25.99142, 24.6487, 24.94563,
    25.2688, 24.41158,
  76.38104, 95.9745, 97.97732, 95.3475, 83.03824, 70.07216, 58.55416,
    54.23248, 45.83961, 42.25657, 48.52514, 47.92913, 50.6848, 50.2244,
    44.24757, 35.54507, 30.07146, 31.52369, 32.9068, 33.94775, 31.36009,
    31.10678, 32.40099, 29.18306, 26.9399, 25.36896, 24.70218, 24.51535,
    24.97005, 24.361,
  56.70181, 64.15337, 60.6856, 56.52192, 49.45416, 52.78687, 70.19624,
    69.60203, 60.00307, 59.60484, 57.32212, 46.15923, 39.06032, 44.47634,
    45.55698, 34.0068, 33.29461, 33.59479, 36.83646, 37.51055, 33.79789,
    31.15856, 28.41878, 25.90338, 25.15445, 25.45169, 24.82539, 24.39217,
    24.41487, 24.13078,
  42.73079, 41.30357, 39.95468, 38.18615, 37.51892, 42.41239, 49.31309,
    47.95965, 44.86864, 43.50868, 41.07887, 34.85267, 31.62774, 35.47927,
    35.10246, 33.06515, 34.15226, 32.72598, 34.17347, 33.46817, 29.14661,
    27.01603, 25.07826, 24.9708, 25.45961, 25.39095, 24.95396, 24.51686,
    24.36347, 24.05979,
  38.95076, 37.16165, 35.80586, 35.41473, 36.4106, 37.12005, 37.27472,
    37.12285, 36.2282, 34.78857, 31.60442, 32.16649, 35.50161, 33.92854,
    32.65685, 32.69905, 32.31973, 30.67863, 32.3789, 30.72502, 25.8837,
    26.20996, 25.72535, 25.09958, 25.14848, 25.39476, 24.88124, 24.29415,
    24.25979, 24.06154,
  35.03623, 34.37822, 33.92918, 34.50109, 34.82075, 35.24472, 35.00702,
    34.64821, 34.02901, 31.58211, 31.72726, 34.9188, 35.40322, 35.04604,
    36.22903, 34.20285, 30.48686, 28.71709, 31.79611, 30.1169, 26.20976,
    26.5721, 26.26256, 25.4976, 24.81391, 25.03353, 24.65417, 24.12593,
    24.08826, 23.97873,
  35.30083, 35.25271, 33.95585, 33.37915, 33.38306, 32.96342, 32.49985,
    32.00021, 30.7794, 29.99481, 32.98033, 33.51266, 30.50093, 31.35259,
    31.94807, 31.1366, 31.10977, 31.91639, 34.55899, 32.89062, 28.9174,
    27.31113, 26.50917, 25.78079, 24.77808, 24.63016, 24.46851, 24.11817,
    24.05841, 23.97642,
  36.00831, 35.73431, 33.90359, 32.3333, 32.1083, 31.63302, 31.08241,
    30.47061, 29.84045, 31.83549, 33.02773, 29.98383, 28.33348, 28.59644,
    28.31603, 27.86983, 29.43212, 31.68161, 33.45814, 33.72245, 31.71319,
    28.75709, 26.72472, 25.99096, 25.16622, 24.64309, 24.41627, 24.14176,
    24.04476, 23.96969,
  35.30752, 35.02924, 33.21951, 31.65355, 31.27497, 31.09008, 30.64862,
    30.01372, 30.07444, 31.99789, 30.4041, 27.31213, 27.89139, 28.26721,
    27.71501, 27.13912, 27.57746, 28.48997, 29.67846, 29.99377, 30.01752,
    29.55022, 28.10213, 26.54886, 25.53723, 24.86583, 24.40018, 24.12515,
    24.06389, 23.9747,
  35.34026, 34.21578, 32.69689, 31.79433, 31.38895, 30.8094, 30.39322,
    29.69345, 30.47707, 30.86626, 27.93968, 26.33132, 27.33767, 27.59987,
    27.32099, 27.07516, 26.75019, 26.76524, 27.11734, 27.14216, 28.14766,
    28.30416, 28.27752, 28.5588, 27.20258, 25.26399, 24.47403, 24.23303,
    24.10116, 23.98927,
  34.92598, 34.14582, 32.32517, 31.49041, 31.88302, 31.9678, 31.28108,
    29.96271, 30.36994, 29.25903, 26.4829, 26.18377, 26.89467, 27.07789,
    26.75708, 27.08887, 26.90084, 26.14787, 26.00059, 26.02433, 26.94181,
    26.82638, 26.49594, 28.12745, 28.49336, 26.08724, 24.72615, 24.64565,
    24.33883, 24.01547,
  34.40042, 33.76916, 32.85068, 32.61084, 32.68064, 32.60922, 32.54742,
    32.08533, 32.22425, 29.22836, 26.37158, 26.81792, 27.51277, 27.93554,
    27.7365, 27.88494, 27.98472, 27.12426, 26.21752, 26.11034, 26.23821,
    26.06357, 25.90244, 26.33272, 27.59716, 27.68641, 26.08086, 24.95759,
    24.69313, 24.12686,
  34.35588, 34.79697, 32.6571, 32.14539, 32.48748, 32.28688, 31.69575,
    31.78434, 32.92697, 29.71006, 26.53296, 27.11146, 27.81123, 28.19583,
    28.46591, 28.58935, 28.23171, 27.82357, 26.86299, 26.08525, 26.13898,
    26.15916, 26.03691, 25.56098, 25.63578, 26.97917, 26.86314, 25.58123,
    25.46007, 24.41013,
  34.66113, 36.52497, 35.13462, 33.57563, 32.38871, 31.48856, 32.21821,
    33.16479, 31.99502, 28.8617, 27.07745, 27.65783, 28.5053, 28.35932,
    28.00994, 28.06239, 27.7721, 27.72917, 27.16751, 26.35867, 26.61495,
    26.63216, 25.72914, 25.22964, 25.32776, 25.92006, 27.15529, 26.22486,
    25.30553, 24.2258,
  35.53098, 37.17471, 34.66286, 33.01818, 32.18447, 31.31359, 32.51717,
    32.80694, 29.94443, 27.66649, 27.46674, 28.06099, 28.48974, 28.16344,
    27.74664, 27.55408, 27.2506, 27.32215, 26.99396, 26.35956, 26.90143,
    27.93407, 27.76807, 26.97018, 26.86842, 26.96185, 28.78683, 28.16793,
    25.23962, 23.84175,
  35.20365, 35.57812, 33.58133, 33.08113, 33.55303, 33.00098, 33.17626,
    31.3162, 28.10452, 27.20733, 27.32822, 27.87759, 28.07937, 27.97468,
    28.10519, 27.80677, 27.14074, 27.05974, 27.46722, 27.73174, 28.47232,
    28.51251, 27.92294, 27.19675, 27.29831, 27.40443, 27.95459, 29.83091,
    27.79587, 24.47052,
  32.86455, 32.18853, 32.70815, 33.86811, 35.16032, 35.96918, 34.10602,
    29.94512, 27.59001, 27.1356, 26.53092, 26.46953, 26.67979, 27.1468,
    27.95208, 28.25973, 28.28493, 28.69494, 28.12577, 27.43493, 27.37777,
    26.9341, 26.17882, 25.80709, 26.13008, 26.63449, 26.69735, 26.74027,
    27.36228, 24.9822,
  32.14961, 32.24082, 32.54731, 32.60995, 33.29994, 35.75498, 35.4422,
    30.37766, 27.51568, 27.60802, 27.92838, 28.42812, 28.97939, 29.30301,
    29.38795, 29.38252, 28.49107, 27.64011, 27.09296, 26.19943, 25.60588,
    25.47849, 25.29015, 25.22366, 25.32249, 25.8779, 25.84227, 25.27394,
    24.99702, 24.16095,
  18.46122, 18.49371, 18.52934, 18.52419, 18.49926, 18.50928, 18.51687,
    18.53985, 18.60678, 18.63697, 19.41404, 19.33362, 18.63773, 18.84473,
    18.89658, 18.63561, 18.57366, 18.59066, 18.59549, 19.10606, 19.26628,
    18.79771, 18.76332, 19.23892, 19.42107, 19.00198, 21.26465, 22.21451,
    20.02979, 19.00712,
  18.79328, 18.73372, 18.63579, 18.81654, 18.65394, 18.55719, 18.60213,
    18.6436, 18.71798, 18.83889, 19.19955, 19.67061, 19.91731, 19.31026,
    19.16823, 19.08935, 18.6951, 18.73341, 19.12902, 19.5654, 19.47799,
    18.88449, 18.89495, 19.5207, 22.901, 22.54647, 22.18099, 24.4893,
    21.05998, 19.60183,
  18.73662, 18.7223, 18.67221, 18.71771, 18.66311, 18.60332, 18.6165,
    18.68196, 18.7693, 18.81504, 18.897, 19.30074, 19.58614, 19.99992,
    19.91639, 19.18302, 19.14705, 19.39989, 19.43493, 19.55007, 20.17407,
    21.10367, 21.91316, 21.29949, 25.86261, 27.34861, 24.0863, 24.2389,
    21.00793, 20.09903,
  18.68398, 18.66863, 18.84387, 18.95789, 19.15481, 19.53325, 19.56608,
    19.35108, 19.38296, 19.58921, 19.59296, 19.92923, 19.73134, 19.51291,
    20.27665, 21.00912, 20.24505, 19.44856, 19.54108, 19.73492, 21.96244,
    22.91243, 22.16702, 26.0762, 26.96376, 25.42105, 26.34651, 23.67006,
    20.83132, 19.50025,
  19.02991, 18.83425, 19.04974, 19.36649, 19.61772, 19.77773, 19.80441,
    19.66522, 20.16537, 20.44999, 20.33947, 20.12049, 19.8506, 20.01603,
    20.61361, 20.99703, 20.02833, 19.49478, 19.8223, 24.10088, 24.80612,
    21.28355, 21.20603, 23.09573, 24.46153, 24.1524, 23.53955, 24.29096,
    24.59757, 20.58473,
  19.04576, 19.10506, 19.79912, 20.74126, 20.57665, 20.10534, 20.24847,
    20.03564, 19.77139, 19.82954, 19.68773, 21.27053, 22.74431, 22.91712,
    22.23744, 28.85065, 33.71196, 26.50616, 22.42364, 24.59125, 22.84748,
    20.11867, 20.61234, 21.20959, 23.76455, 22.98962, 26.24896, 36.81157,
    32.22152, 20.16049,
  19.1898, 19.49501, 20.30483, 21.15709, 21.13481, 20.71689, 21.52817,
    22.86802, 23.07393, 23.06164, 23.50935, 23.09859, 22.4132, 22.49728,
    27.20535, 33.48501, 31.24138, 24.41515, 22.37174, 22.14749, 20.86688,
    20.11846, 20.57652, 22.69054, 24.08636, 21.79832, 31.50277, 44.2994,
    32.41159, 19.0254,
  19.4556, 19.79202, 20.74397, 21.56935, 21.38082, 23.29144, 25.24388,
    23.56644, 22.49045, 22.61053, 22.58777, 21.65166, 20.90231, 21.00859,
    23.48528, 24.91975, 23.56204, 22.06431, 21.02094, 20.83927, 20.35198,
    20.17052, 21.32239, 23.57813, 23.38595, 21.60733, 34.58179, 38.09933,
    24.40657, 19.18917,
  21.05832, 21.28989, 22.45935, 22.5675, 23.09431, 24.9407, 24.05451,
    22.45551, 22.51657, 22.63166, 22.05042, 21.19438, 20.74219, 23.92373,
    24.93759, 22.20474, 22.41132, 23.60256, 23.57938, 21.63948, 20.25104,
    21.42718, 25.30639, 25.80832, 23.08158, 23.15193, 29.75217, 27.94046,
    20.99433, 19.23918,
  23.69455, 25.05036, 26.91261, 28.05535, 28.2992, 25.13581, 21.87826,
    21.66061, 21.58479, 21.0298, 22.21887, 25.0272, 26.25298, 26.01552,
    24.97395, 24.82499, 25.4196, 25.92906, 24.97034, 23.98409, 23.93771,
    24.8832, 26.08469, 24.71135, 29.5021, 36.84914, 30.57721, 22.03932,
    19.78433, 18.69391,
  34.12499, 36.53513, 33.88528, 29.54443, 29.01081, 27.58994, 24.50274,
    25.90356, 27.40904, 34.14831, 35.56868, 26.12569, 23.86141, 23.42635,
    22.90956, 23.85763, 25.02033, 25.13776, 24.17103, 24.41828, 26.79386,
    26.74066, 23.81574, 21.91565, 26.00656, 29.80095, 24.21029, 19.48987,
    18.982, 18.57296,
  45.52654, 36.79146, 38.6534, 40.01128, 38.29951, 34.53458, 36.38042,
    33.11789, 28.52479, 33.17123, 31.71598, 22.15399, 23.12343, 23.98003,
    22.99487, 23.3545, 23.06332, 23.10731, 22.81413, 23.5883, 26.72898,
    25.51609, 21.60506, 24.78812, 26.06013, 21.16369, 19.03531, 19.28922,
    19.23064, 18.71546,
  51.18813, 50.22982, 66.57664, 71.16718, 69.73058, 61.01066, 45.53868,
    31.75564, 29.38521, 27.93594, 24.65969, 20.80387, 25.14496, 26.97851,
    24.15247, 23.51166, 23.55932, 22.96979, 22.64442, 25.07503, 26.76773,
    24.02571, 21.31251, 26.42082, 26.98446, 20.54808, 19.18113, 19.49567,
    19.78309, 18.96488,
  62.59727, 86.32122, 86.86099, 80.34009, 69.68228, 60.37889, 52.21223,
    45.77937, 36.93214, 34.16746, 39.3921, 39.6285, 43.30075, 43.21455,
    36.73748, 28.41977, 24.12428, 25.55678, 27.04765, 28.1477, 25.70783,
    25.47696, 26.74758, 23.88399, 21.56562, 19.85405, 19.26821, 19.09154,
    19.52757, 18.94211,
  48.71639, 57.17918, 54.80807, 50.77725, 43.61306, 47.68288, 63.47828,
    61.1736, 51.45267, 51.77384, 50.52285, 39.74845, 33.35485, 38.78221,
    38.71429, 27.83788, 27.17397, 27.25353, 29.55494, 30.56558, 28.16537,
    25.84708, 23.4376, 20.66908, 19.60603, 19.90909, 19.33079, 18.94586,
    18.99445, 18.71479,
  36.34785, 36.17082, 35.60457, 34.22582, 32.9904, 38.32687, 45.53151,
    42.9505, 39.98692, 39.33125, 36.00911, 28.86343, 25.31528, 29.60809,
    29.33851, 27.04712, 28.28833, 26.53199, 27.31621, 27.07744, 23.92452,
    21.81825, 19.77144, 19.67319, 20.01164, 19.8396, 19.44393, 19.05926,
    18.93457, 18.65386,
  33.59519, 32.43184, 31.1488, 30.5668, 31.18936, 31.82026, 31.9765,
    31.31209, 30.40046, 28.97105, 25.521, 26.02763, 28.84887, 27.60322,
    26.95741, 27.04877, 26.80964, 24.78465, 25.76482, 24.43418, 20.41495,
    20.67953, 20.26791, 19.78603, 19.76317, 19.85871, 19.37282, 18.8675,
    18.84256, 18.63986,
  30.27863, 29.50984, 28.76034, 29.25812, 29.74818, 30.41099, 30.39339,
    29.90384, 28.77074, 26.02649, 25.49186, 28.6817, 29.77141, 29.26882,
    30.51245, 28.79602, 25.11726, 23.04618, 25.38334, 23.79614, 20.51163,
    20.79576, 20.57118, 20.04432, 19.43793, 19.56331, 19.18733, 18.7007,
    18.67882, 18.57766,
  30.00089, 29.98415, 28.86324, 28.73788, 29.13402, 29.15491, 28.82806,
    27.87758, 25.9632, 24.51463, 26.98598, 27.86493, 25.50411, 26.28943,
    26.83381, 25.98842, 25.51683, 25.76831, 27.55077, 25.81617, 22.74191,
    21.42242, 20.68667, 20.20227, 19.36548, 19.2304, 19.03711, 18.69307,
    18.64963, 18.56258,
  30.79546, 30.97385, 29.49064, 28.39027, 28.5129, 28.16422, 27.47146,
    26.36753, 24.98092, 26.26484, 27.38315, 24.77441, 23.17332, 23.24276,
    22.92001, 22.56467, 23.89326, 25.75564, 26.71712, 26.62457, 25.32318,
    22.79443, 20.85852, 20.37117, 19.67798, 19.2076, 18.98635, 18.726,
    18.65445, 18.56493,
  30.64088, 30.99943, 29.46255, 28.12057, 27.85705, 27.62392, 27.01593,
    26.0208, 25.43184, 26.84673, 25.30179, 22.23223, 22.62583, 22.65628,
    21.99134, 21.54558, 21.96199, 22.77202, 23.45263, 23.63979, 24.10435,
    23.71298, 22.20358, 20.92826, 20.05814, 19.40513, 18.99141, 18.72706,
    18.65126, 18.56288,
  31.12783, 30.64588, 29.12484, 28.26007, 27.90149, 27.37507, 26.9709,
    26.05174, 26.06101, 26.00614, 23.02523, 21.0243, 21.80758, 21.90262,
    21.55855, 21.4146, 21.17379, 21.10771, 21.42288, 21.51143, 22.49672,
    22.52182, 22.31787, 22.51018, 21.31012, 19.70173, 19.04153, 18.81144,
    18.68137, 18.57212,
  31.04035, 30.62832, 28.77019, 27.98227, 28.45699, 28.63033, 28.01988,
    26.39394, 25.97968, 24.48985, 21.45671, 20.66894, 21.24777, 21.38144,
    21.1038, 21.47541, 21.30687, 20.59462, 20.50476, 20.50731, 21.46119,
    21.2142, 20.72167, 22.25101, 22.5456, 20.42592, 19.28165, 19.21777,
    18.9096, 18.60074,
  30.48354, 30.2393, 29.31127, 29.19394, 29.47843, 29.56745, 29.38959,
    28.50518, 27.6747, 24.0735, 21.05725, 21.19831, 21.83181, 22.18777,
    21.97282, 22.16463, 22.23604, 21.36042, 20.63132, 20.65457, 20.73954,
    20.45964, 20.2324, 20.67752, 21.83479, 22.11129, 20.66092, 19.55195,
    19.27286, 18.70362,
  30.63232, 31.34194, 29.48846, 29.01332, 29.44494, 29.32918, 28.67873,
    28.10673, 28.18737, 24.45943, 21.14025, 21.49817, 22.09743, 22.46864,
    22.6813, 22.74187, 22.36918, 21.93154, 21.22518, 20.68439, 20.55772,
    20.51536, 20.45329, 20.06398, 20.23483, 21.74899, 21.60625, 20.24665,
    20.06795, 18.99396,
  31.13731, 33.27262, 31.73215, 30.07009, 29.18093, 28.37092, 28.91458,
    29.29202, 27.29123, 23.76119, 21.68814, 21.92756, 22.57706, 22.52785,
    22.26755, 22.27939, 21.89706, 21.81439, 21.49718, 20.90719, 20.96705,
    20.94448, 20.19756, 19.78081, 19.90818, 20.6403, 21.81771, 20.80228,
    19.95728, 18.86961,
  32.26643, 34.2882, 31.62062, 29.6167, 28.70565, 28.00388, 29.4251,
    29.21885, 25.45152, 22.6412, 22.08606, 22.31609, 22.61617, 22.37757,
    21.99326, 21.80045, 21.45624, 21.48638, 21.34731, 20.89762, 21.18944,
    22.04131, 21.85384, 21.30145, 21.36871, 21.56287, 23.47044, 22.67629,
    19.81292, 18.48341,
  32.10688, 32.78782, 30.20289, 29.21426, 29.67036, 29.3453, 29.61941,
    27.48379, 23.64568, 22.11288, 21.95005, 22.17484, 22.23643, 22.19212,
    22.27516, 21.93623, 21.33215, 21.21286, 21.79698, 22.31751, 22.66837,
    22.5661, 22.095, 21.64909, 21.89457, 21.99602, 22.6864, 24.43356,
    22.26958, 19.03287,
  29.70494, 28.98115, 29.31999, 30.52916, 31.45592, 31.84408, 30.28963,
    26.04222, 22.97531, 21.90898, 21.10298, 20.94923, 21.11222, 21.40041,
    21.93494, 22.13972, 22.16453, 22.53518, 22.4396, 22.15884, 22.0211,
    21.52139, 20.73846, 20.40652, 20.74627, 21.23199, 21.2694, 21.40848,
    22.01918, 19.55062,
  28.56552, 28.70304, 29.194, 29.49504, 30.06699, 31.79235, 30.96268,
    25.94325, 22.61015, 22.08657, 22.07369, 22.58235, 23.13667, 23.07989,
    23.03224, 23.16236, 22.41888, 21.76071, 21.50915, 20.81019, 20.27067,
    20.1274, 19.8831, 19.79578, 19.90849, 20.46362, 20.48421, 19.85838,
    19.60577, 18.78104,
  15.57024, 15.59912, 15.62722, 15.61657, 15.61231, 15.60798, 15.60487,
    15.62358, 15.68625, 15.69851, 16.42619, 16.30783, 15.70876, 15.90378,
    15.94433, 15.71779, 15.66771, 15.68444, 15.66538, 16.11043, 16.19358,
    15.79149, 15.78072, 16.19575, 16.29381, 15.88631, 18.04755, 18.70371,
    16.93145, 16.06913,
  15.87987, 15.7998, 15.73174, 15.86969, 15.73079, 15.64726, 15.6724,
    15.70804, 15.78409, 15.90154, 16.36355, 16.74438, 16.8857, 16.3276,
    16.27027, 16.13725, 15.77223, 15.79431, 16.15364, 16.56924, 16.47307,
    15.88047, 15.85985, 16.42463, 19.49121, 18.76523, 19.29652, 21.29049,
    18.06388, 16.64592,
  15.87261, 15.8274, 15.76777, 15.82018, 15.74565, 15.67044, 15.68753,
    15.7505, 15.85071, 15.90946, 15.97437, 16.40474, 16.70994, 17.02295,
    16.90344, 16.20703, 16.12555, 16.32256, 16.40315, 16.46432, 16.94502,
    17.71559, 18.48895, 17.8285, 22.43517, 23.45431, 21.01979, 21.11643,
    18.05456, 17.11441,
  15.7505, 15.74745, 15.88975, 15.96887, 16.16615, 16.48757, 16.50164,
    16.3294, 16.35562, 16.4964, 16.49704, 16.91053, 16.67919, 16.58171,
    17.22122, 17.77874, 17.01505, 16.31686, 16.33019, 16.3651, 18.54364,
    19.46194, 18.96359, 22.57987, 23.26593, 22.60864, 23.42535, 20.50691,
    17.75909, 16.57131,
  16.00599, 15.87007, 16.04118, 16.34707, 16.57371, 16.76981, 16.80249,
    16.59742, 17.08329, 17.37038, 17.28962, 17.04262, 16.76751, 16.87117,
    17.42912, 17.80546, 16.63515, 16.09955, 16.40925, 20.21276, 20.85411,
    18.22885, 18.1306, 20.36272, 21.4702, 21.1233, 20.69202, 21.03917,
    20.94091, 17.3439,
  16.01623, 16.02396, 16.66668, 17.52975, 17.4192, 17.00043, 17.12257,
    16.92946, 16.73989, 16.80104, 16.50613, 17.91592, 19.2062, 19.38101,
    18.52648, 23.9704, 27.71313, 21.8838, 18.75431, 21.23945, 19.5528,
    17.12549, 17.68306, 18.13516, 20.77553, 19.77206, 22.45768, 31.79568,
    27.66764, 17.10468,
  16.07011, 16.33293, 17.15271, 17.9846, 18.02505, 17.42068, 18.07523,
    19.25529, 19.27716, 19.23666, 19.63721, 19.44778, 18.99271, 18.96668,
    23.05722, 28.80945, 27.41032, 21.16143, 19.20106, 19.05502, 17.81328,
    17.12365, 17.57788, 19.57837, 20.89741, 18.41088, 27.86987, 39.90178,
    28.45451, 16.08983,
  16.24334, 16.52891, 17.4328, 18.18806, 17.95692, 19.49774, 21.12383,
    19.80146, 18.98254, 19.08891, 19.23721, 18.21286, 17.44856, 17.45825,
    20.39501, 21.97247, 20.46113, 18.84954, 17.96708, 17.82388, 17.35806,
    17.16349, 18.11202, 20.30902, 20.13554, 18.1346, 31.44309, 34.57035,
    21.43641, 16.19894,
  17.29727, 17.45955, 18.50924, 18.4639, 18.93329, 20.97987, 20.3325,
    18.77441, 18.84173, 18.92704, 18.36339, 17.58194, 17.19124, 20.42527,
    21.33019, 18.94021, 19.33916, 20.36789, 20.16385, 18.33334, 17.12609,
    18.11339, 21.65513, 22.00811, 19.6976, 19.55981, 26.95133, 24.81105,
    17.98679, 16.30212,
  19.04859, 20.13358, 22.07585, 23.06919, 23.46892, 20.59542, 17.94704,
    17.85003, 18.06303, 17.44918, 18.59356, 21.1734, 22.36066, 22.52639,
    21.88628, 21.56409, 21.92005, 22.37604, 21.65855, 20.76081, 20.49433,
    21.44828, 22.82608, 21.57341, 25.763, 32.41504, 27.02536, 19.30746,
    16.96251, 15.81513,
  27.00194, 29.44926, 27.73772, 24.05353, 24.03944, 22.3552, 19.71257,
    21.45245, 22.60331, 29.17035, 30.47846, 22.93316, 20.99519, 20.41253,
    19.79302, 20.83219, 22.00247, 22.01282, 20.93905, 21.34011, 23.63142,
    23.6169, 20.75348, 19.06466, 23.49225, 27.74227, 21.80408, 16.72299,
    16.07475, 15.67401,
  36.94072, 30.49446, 31.00373, 31.4581, 29.78246, 27.12954, 29.35671,
    27.52254, 24.30346, 29.62137, 28.39662, 19.42716, 19.9614, 20.75528,
    20.03193, 20.31, 20.05768, 20.11314, 19.71797, 20.49216, 23.81293,
    22.53924, 18.74105, 21.73661, 22.8837, 18.43689, 16.23993, 16.38392,
    16.31044, 15.8092,
  46.03087, 41.9128, 49.76085, 55.43117, 55.49085, 49.94825, 37.99926,
    26.8019, 25.3455, 24.45278, 21.08819, 17.71788, 21.87872, 23.60034,
    21.13863, 20.48229, 20.55945, 19.90858, 19.57502, 22.08255, 23.94566,
    21.1896, 18.4146, 23.80233, 24.07079, 17.71765, 16.2706, 16.61749,
    16.89095, 16.04286,
  55.30519, 72.06281, 74.08828, 73.60574, 69.82539, 58.39313, 43.3918,
    38.67307, 30.64205, 28.72486, 33.07998, 33.86716, 38.10347, 38.68745,
    32.92348, 25.14915, 21.26266, 22.57788, 23.99271, 25.14646, 22.84255,
    22.52486, 23.51239, 21.25368, 18.92777, 16.95967, 16.34369, 16.22013,
    16.71821, 16.03402,
  41.6664, 50.01711, 50.59211, 49.63913, 44.01621, 43.80799, 53.88535,
    52.20272, 42.23511, 43.80866, 44.34563, 35.4487, 30.45182, 35.62122,
    34.95983, 25.20235, 24.32787, 24.24734, 26.33696, 27.27114, 25.0623,
    23.08723, 20.95485, 17.93001, 16.70802, 17.01171, 16.42459, 16.03588,
    16.13576, 15.81882,
  29.38527, 30.14309, 30.65597, 29.5704, 27.30989, 32.47137, 39.8674,
    36.74017, 34.43484, 35.25653, 32.67809, 25.62472, 22.26379, 26.66776,
    26.31519, 24.34622, 25.69437, 23.62683, 24.31568, 24.24443, 21.48941,
    19.17263, 16.94098, 16.83026, 17.12818, 16.89881, 16.54791, 16.16077,
    16.02556, 15.75104,
  27.85907, 27.15732, 25.9475, 24.96038, 25.19911, 25.95285, 26.41691,
    25.90497, 25.86961, 25.2304, 22.20757, 22.84075, 25.28101, 24.29268,
    24.01262, 24.35402, 24.35328, 22.03197, 23.00962, 21.51777, 17.62354,
    17.7895, 17.37964, 16.90733, 16.85873, 16.92165, 16.46266, 15.97987,
    15.95226, 15.73691,
  25.11905, 24.19749, 23.24096, 23.5181, 23.95387, 24.56086, 24.92522,
    24.99735, 24.33258, 22.19617, 21.76584, 25.09736, 26.38534, 26.10193,
    27.74977, 26.20072, 22.51643, 20.20784, 22.56008, 20.72724, 17.53823,
    17.78248, 17.60759, 17.02842, 16.48219, 16.67045, 16.26855, 15.79274,
    15.77684, 15.67763,
  24.52484, 24.14922, 22.92352, 22.78453, 23.2184, 23.47865, 23.48131,
    22.95455, 21.54348, 20.61286, 23.33813, 24.46079, 22.73732, 23.8129,
    24.38988, 23.40458, 22.50867, 22.32132, 24.17403, 22.39711, 19.53889,
    18.25432, 17.60019, 17.1238, 16.36584, 16.32825, 16.12748, 15.77568,
    15.73731, 15.66054,
  25.0942, 24.9552, 23.41356, 22.45351, 22.67274, 22.43193, 22.04011,
    21.43043, 20.65977, 22.43921, 23.85505, 21.79587, 20.45884, 20.52377,
    20.12282, 19.67853, 20.97549, 22.6978, 23.6909, 23.74947, 22.3546,
    19.61074, 17.6763, 17.26022, 16.67412, 16.25147, 16.06572, 15.80024,
    15.73027, 15.65737,
  24.7715, 24.97288, 23.43521, 22.25137, 22.12013, 21.98955, 21.64568,
    21.17633, 21.27171, 23.46371, 22.27562, 19.58219, 19.89493, 19.73201,
    19.01771, 18.56149, 19.03742, 19.88799, 20.60379, 20.93222, 21.59837,
    20.67894, 18.81066, 17.77527, 17.03903, 16.40721, 16.05927, 15.81879,
    15.73767, 15.65168,
  25.10524, 24.61814, 23.22486, 22.47721, 22.18767, 21.86056, 21.74517,
    21.42857, 22.13733, 22.83465, 20.22824, 18.25286, 18.88714, 18.92117,
    18.55794, 18.43137, 18.24534, 18.23417, 18.63278, 18.71733, 19.7673,
    19.52484, 19.24193, 19.25384, 18.10785, 16.67265, 16.10111, 15.86921,
    15.7639, 15.66207,
  25.17323, 24.6935, 23.01877, 22.38133, 22.84444, 23.16217, 22.90531,
    21.86056, 22.17715, 21.35426, 18.63682, 17.74131, 18.22803, 18.32364,
    18.1024, 18.46133, 18.27726, 17.66007, 17.66948, 17.6914, 18.58605,
    18.11693, 17.76971, 19.18524, 19.30776, 17.30636, 16.34516, 16.26936,
    15.97113, 15.68207,
  24.79966, 24.58879, 23.58807, 23.50573, 23.95329, 24.32324, 24.44226,
    24.02531, 23.65135, 20.56552, 18.02252, 18.1062, 18.67545, 19.04366,
    18.84366, 18.97409, 19.01796, 18.20861, 17.62943, 17.71075, 17.80531,
    17.47231, 17.19756, 17.66649, 18.78469, 18.8809, 17.51242, 16.61426,
    16.30025, 15.76082,
  25.00072, 25.26014, 23.82007, 23.67135, 24.28114, 24.48336, 24.08903,
    23.72883, 24.09122, 20.7911, 18.02515, 18.4177, 19.00846, 19.36616,
    19.54978, 19.47568, 19.16467, 18.81656, 18.18563, 17.75028, 17.62152,
    17.49786, 17.47305, 17.093, 17.32898, 18.86029, 18.60908, 17.25162,
    17.13215, 16.0262,
  25.46352, 27.02724, 25.89289, 24.70069, 24.09395, 23.49236, 23.93822,
    24.25302, 22.89144, 20.14553, 18.44651, 18.84397, 19.48129, 19.37845,
    19.17389, 19.12975, 18.72625, 18.74531, 18.47848, 17.94055, 17.99949,
    17.96369, 17.25119, 16.90803, 16.99634, 17.78391, 19.01677, 17.79639,
    17.10878, 15.94657,
  26.76574, 28.42176, 26.43225, 24.70391, 23.50147, 22.68159, 24.14052,
    24.22866, 21.20093, 19.16794, 18.89491, 19.28577, 19.57604, 19.26036,
    18.88601, 18.69971, 18.36917, 18.45251, 18.34855, 17.9305, 18.14849,
    18.99715, 18.69646, 18.2712, 18.37203, 18.48416, 20.60538, 19.57408,
    16.8079, 15.57427,
  27.26813, 27.75585, 25.03186, 23.94709, 24.0192, 23.63897, 24.15742,
    22.58821, 19.64129, 18.72862, 18.86729, 19.15344, 19.17977, 19.10769,
    19.21103, 18.85003, 18.25814, 18.16937, 18.764, 19.19127, 19.47309,
    19.44997, 19.0741, 18.66994, 18.97163, 18.95115, 19.82988, 21.63181,
    19.21419, 16.0603,
  25.03872, 23.92169, 23.96899, 24.96291, 25.58071, 25.7997, 24.787,
    21.32116, 19.14748, 18.61539, 18.08674, 17.97901, 18.07738, 18.35995,
    18.9392, 19.09304, 19.02102, 19.33163, 19.33126, 19.17816, 19.08671,
    18.5614, 17.78671, 17.47536, 17.85242, 18.33101, 18.38024, 18.87256,
    19.43945, 16.56951,
  23.59495, 23.26418, 23.82066, 24.19194, 24.64278, 26.09873, 25.449,
    21.29571, 18.87835, 18.72926, 18.79097, 19.18213, 19.62722, 19.63124,
    19.68252, 19.92646, 19.24239, 18.71745, 18.51784, 17.8269, 17.35859,
    17.26729, 16.97691, 16.88805, 17.01223, 17.6168, 17.66385, 17.06401,
    16.91839, 15.9069,
  14.07755, 14.10796, 14.12765, 14.12942, 14.12629, 14.13251, 14.12317,
    14.13068, 14.18174, 14.18699, 14.89343, 14.84035, 14.21166, 14.38568,
    14.4644, 14.2514, 14.20165, 14.19616, 14.15635, 14.59285, 14.74084,
    14.3613, 14.32764, 14.71784, 14.79349, 14.38858, 16.53809, 17.41059,
    15.54789, 14.64877,
  14.32981, 14.29562, 14.23146, 14.39868, 14.26154, 14.17062, 14.19153,
    14.21732, 14.2859, 14.40831, 14.9829, 15.38702, 15.43473, 14.91214,
    14.81153, 14.70963, 14.32149, 14.30262, 14.65787, 15.1858, 15.14326,
    14.46201, 14.35185, 14.91384, 17.9686, 17.6141, 18.08931, 20.60815,
    16.87933, 15.31315,
  14.3817, 14.36221, 14.30877, 14.3928, 14.29018, 14.17956, 14.18734,
    14.26413, 14.36448, 14.45061, 14.53581, 15.0044, 15.39002, 15.63337,
    15.49967, 14.77481, 14.64326, 14.87432, 14.9731, 15.04451, 15.4054,
    16.08678, 16.78679, 16.15495, 20.96119, 22.82257, 20.1218, 20.57266,
    16.87724, 15.83579,
  14.26379, 14.26904, 14.41026, 14.45547, 14.64108, 14.97808, 14.97606,
    14.80501, 14.83016, 14.98679, 15.07261, 15.50674, 15.24891, 15.17734,
    15.84205, 16.35461, 15.6766, 14.88504, 14.78049, 14.68863, 16.89742,
    18.02708, 17.43548, 21.119, 22.45624, 21.91539, 23.134, 20.0649,
    16.65339, 15.289,
  14.55653, 14.36766, 14.52267, 14.78593, 15.05491, 15.36202, 15.3649,
    15.11108, 15.61426, 16.0396, 16.02973, 15.73008, 15.29472, 15.38372,
    16.07101, 16.53291, 15.24055, 14.39506, 14.61884, 18.48646, 19.6868,
    16.85992, 16.6666, 19.40536, 20.69881, 20.30223, 20.22213, 20.27935,
    19.95251, 16.11518,
  14.55598, 14.46241, 15.03348, 15.91606, 15.99825, 15.63705, 15.65184,
    15.48485, 15.38383, 15.47918, 15.17331, 16.46928, 17.79883, 17.94879,
    17.05466, 21.80667, 25.72029, 20.27881, 17.10438, 20.15477, 18.6692,
    15.67135, 16.33896, 16.9729, 19.80322, 19.02026, 20.84823, 30.74906,
    27.60131, 15.91695,
  14.49136, 14.72579, 15.57838, 16.53887, 16.72327, 16.09189, 16.55789,
    17.817, 17.77638, 17.69646, 18.15647, 18.18491, 17.77127, 17.51666,
    21.22759, 27.64504, 26.90686, 20.17478, 18.00096, 17.98693, 16.59488,
    15.7799, 16.29045, 18.48403, 20.001, 17.40915, 26.16891, 39.94175,
    29.15541, 14.71874,
  14.64163, 14.96779, 15.94426, 16.78248, 16.5407, 17.8294, 19.62067,
    18.6013, 17.77012, 17.90602, 18.13053, 16.95765, 15.81363, 15.68092,
    18.97793, 21.32998, 19.65799, 17.7062, 16.74837, 16.55777, 16.08686,
    15.85105, 16.81801, 19.3345, 19.16467, 16.9516, 30.73849, 35.64364,
    21.10711, 14.78432,
  15.6755, 15.85996, 17.01143, 16.98356, 17.32768, 19.65454, 19.23722,
    17.416, 17.47388, 17.63114, 16.94079, 15.89816, 15.30596, 18.63544,
    20.10201, 17.71998, 18.15427, 19.47367, 19.27107, 17.22859, 15.74451,
    16.76905, 20.51558, 21.16346, 18.5756, 18.43266, 26.71454, 24.90711,
    16.66476, 14.92634,
  17.70748, 18.62357, 20.63333, 21.85755, 22.27413, 19.5196, 16.58744,
    16.40212, 16.63411, 15.90984, 16.84529, 19.56088, 20.97195, 21.43833,
    20.94103, 20.48112, 20.91248, 21.68053, 21.07738, 19.80184, 19.23714,
    20.26598, 21.9612, 20.70118, 24.23235, 31.42707, 26.76586, 18.35274,
    15.65713, 14.37996,
  23.40352, 26.48216, 26.28284, 23.09796, 23.10173, 21.38388, 18.41992,
    20.04734, 20.88298, 26.78764, 28.84339, 21.90273, 20.14197, 19.45416,
    18.63911, 19.89979, 21.26888, 21.37152, 20.17022, 20.33257, 22.8077,
    22.75358, 19.70675, 17.88407, 22.58429, 27.60016, 21.5373, 15.46585,
    14.6406, 14.18169,
  37.66751, 30.76903, 28.28417, 29.3041, 27.52558, 24.56549, 27.05576,
    26.00688, 22.76704, 28.16417, 27.73569, 18.26396, 18.61925, 19.59967,
    19.03448, 19.41448, 19.09593, 19.10547, 18.72263, 19.5318, 23.0254,
    21.65864, 17.47147, 20.46203, 22.14067, 17.52738, 14.88484, 14.93043,
    14.83999, 14.3275,
  50.33471, 39.54741, 43.89178, 50.71008, 50.72551, 46.14458, 35.93591,
    25.1962, 24.1439, 23.59066, 20.21907, 16.2131, 20.57742, 22.5811,
    20.1088, 19.42178, 19.44506, 18.73333, 18.52915, 21.41915, 23.40654,
    20.14808, 17.19042, 22.98238, 23.83382, 16.6108, 14.81521, 15.20029,
    15.39474, 14.57015,
  54.91169, 65.78798, 67.66899, 69.1516, 65.32435, 55.10917, 41.82452,
    37.48756, 29.80676, 27.20137, 31.76174, 32.17097, 36.2985, 36.99781,
    31.77819, 24.28762, 20.16668, 21.55418, 23.395, 24.94821, 22.47447,
    21.3909, 22.68592, 20.78876, 18.20303, 15.63647, 14.92624, 14.82656,
    15.2788, 14.59379,
  38.81297, 45.98293, 47.40425, 48.42143, 43.27288, 41.32753, 50.88597,
    50.52978, 40.37152, 42.03721, 43.37352, 34.76289, 29.61314, 34.7373,
    34.76348, 24.47064, 23.488, 23.57846, 25.97569, 27.15829, 24.58027,
    22.47376, 20.57065, 17.11716, 15.27059, 15.62646, 15.01493, 14.61852,
    14.72776, 14.38278,
  25.93207, 26.98544, 28.4485, 28.12207, 25.59963, 30.21285, 37.87951,
    34.83235, 32.83153, 34.63822, 32.45678, 25.01398, 21.31304, 26.1174,
    25.99477, 23.73966, 25.28427, 23.16445, 23.83188, 24.07353, 21.05887,
    18.53347, 15.97936, 15.64612, 15.78991, 15.50409, 15.13471, 14.76979,
    14.60233, 14.29012,
  24.76477, 24.40837, 23.5048, 22.20806, 22.13281, 23.54258, 24.61384,
    24.02112, 24.42226, 24.42648, 21.38731, 21.9539, 24.63678, 23.40163,
    23.27618, 23.97331, 24.11338, 21.61854, 22.47448, 21.28367, 16.65259,
    16.55609, 16.16636, 15.7478, 15.54311, 15.50227, 15.05808, 14.5808,
    14.53116, 14.28708,
  22.26171, 21.42951, 20.34093, 20.5005, 21.06493, 21.9237, 22.64846,
    23.11565, 22.80059, 20.81036, 20.32445, 24.37806, 25.99047, 25.18113,
    27.41546, 26.01398, 22.17282, 19.4687, 21.98126, 20.3159, 16.25895,
    16.47847, 16.33745, 15.81573, 15.13703, 15.25843, 14.87633, 14.34587,
    14.33245, 14.21905,
  21.76257, 21.23807, 19.9132, 19.78098, 20.27833, 20.78878, 21.10788,
    20.92484, 19.85133, 19.00123, 22.05058, 23.80942, 21.97238, 23.22533,
    24.55964, 23.54996, 22.04655, 21.30193, 23.47046, 21.57722, 18.12839,
    16.91081, 16.2772, 15.8157, 14.97641, 14.89822, 14.70297, 14.31996,
    14.26463, 14.18456,
  22.30983, 21.99341, 20.39369, 19.40379, 19.70591, 19.67539, 19.54651,
    19.23825, 18.7272, 20.83588, 22.9515, 21.04418, 19.5169, 19.95714,
    19.93843, 19.5262, 20.61755, 22.01828, 22.98189, 22.97746, 21.18953,
    18.40221, 16.37617, 15.92874, 15.29202, 14.82013, 14.61757, 14.35715,
    14.26599, 14.18077,
  21.81205, 21.92814, 20.43665, 19.26204, 19.20493, 19.1815, 18.99225,
    18.84109, 19.42764, 22.34206, 21.73611, 18.82205, 19.12825, 19.07249,
    18.34938, 17.76367, 18.19654, 18.92909, 19.6785, 20.17837, 20.79402,
    19.737, 17.57463, 16.52022, 15.72896, 15.02664, 14.6262, 14.35545,
    14.27321, 14.18794,
  22.15808, 21.57882, 20.28052, 19.54016, 19.23969, 18.92093, 19.04476,
    19.29179, 20.6969, 22.12598, 19.74845, 17.53658, 18.153, 18.06625,
    17.53353, 17.24143, 17.05296, 17.13126, 17.63767, 17.67656, 18.86778,
    18.73344, 18.18894, 18.27225, 16.97088, 15.34077, 14.6709, 14.42171,
    14.28582, 14.18269,
  22.36667, 21.71712, 20.10743, 19.42902, 19.86559, 20.3357, 20.45413,
    19.9759, 21.12791, 20.9138, 18.05749, 16.92118, 17.30572, 17.24284,
    16.91491, 17.29784, 17.2572, 16.65885, 16.53854, 16.48434, 17.59146,
    17.17839, 16.65314, 18.29918, 18.34547, 16.05999, 14.90391, 14.82609,
    14.52192, 14.21144,
  22.12623, 21.66854, 20.58194, 20.53719, 21.14898, 21.84377, 22.58593,
    22.72846, 22.84913, 19.96214, 17.10224, 17.01136, 17.54268, 17.93873,
    17.73219, 17.95947, 18.13599, 17.19156, 16.35603, 16.4302, 16.68353,
    16.31808, 15.90729, 16.50178, 17.73381, 17.63542, 16.12929, 15.22968,
    14.8871, 14.30126,
  22.18534, 22.07408, 20.82346, 20.97653, 22.03247, 22.62381, 22.66178,
    22.77765, 23.33138, 19.96372, 16.86322, 17.25744, 17.95656, 18.45827,
    18.61583, 18.51047, 18.23592, 17.82597, 17.00711, 16.48607, 16.3088,
    16.18516, 16.19746, 15.78475, 16.05625, 17.65686, 17.39154, 15.92539,
    15.73395, 14.62248,
  22.38785, 23.50596, 22.92394, 22.38563, 22.25618, 22.02913, 22.53796,
    23.04259, 21.9108, 19.18406, 17.19731, 17.69613, 18.50733, 18.44905,
    18.16109, 18.05759, 17.66793, 17.67442, 17.33509, 16.65841, 16.64169,
    16.63283, 15.97041, 15.55606, 15.59368, 16.46704, 17.79988, 16.55654,
    15.77442, 14.58748,
  23.58813, 24.91557, 23.96229, 22.82562, 21.66918, 20.86672, 22.69369,
    23.20062, 20.10254, 18.01029, 17.74976, 18.21861, 18.63142, 18.22603,
    17.70915, 17.53444, 17.22784, 17.28822, 17.10638, 16.61937, 16.84307,
    17.73405, 17.48461, 16.9596, 17.04932, 17.21215, 19.35418, 18.35484,
    15.48873, 14.17371,
  24.93287, 25.20025, 22.70309, 22.01153, 21.96783, 21.65025, 22.54597,
    21.35039, 18.33806, 17.52679, 17.75359, 18.05853, 18.06431, 17.89435,
    17.95786, 17.6371, 16.99144, 16.87551, 17.44452, 17.91341, 18.29577,
    18.37732, 17.97639, 17.51134, 17.82529, 17.79819, 18.67447, 20.5149,
    18.12157, 14.70237,
  23.35595, 22.0505, 21.82513, 22.95181, 23.54636, 23.79024, 22.98014,
    19.82734, 17.83969, 17.54706, 16.97659, 16.77224, 16.82214, 17.13316,
    17.741, 17.84066, 17.6832, 18.00902, 18.09441, 18.03897, 18.03184,
    17.46285, 16.57245, 16.21159, 16.63029, 17.07705, 17.13689, 17.74482,
    18.36411, 15.28983,
  21.81558, 21.23489, 21.72795, 22.14136, 22.59874, 24.17197, 23.71231,
    19.84959, 17.64913, 17.66293, 17.61127, 17.87933, 18.34937, 18.48756,
    18.55637, 18.71733, 18.03785, 17.52936, 17.319, 16.59282, 16.10614,
    15.98664, 15.63948, 15.50427, 15.65075, 16.27729, 16.37299, 15.71815,
    15.59161, 14.51655,
  17.64818, 17.67759, 17.68055, 17.68461, 17.68019, 17.67369, 17.67265,
    17.70209, 17.74063, 17.75274, 18.46281, 18.51735, 17.80146, 17.95715,
    18.06559, 17.84439, 17.7864, 17.78224, 17.74279, 18.13836, 18.33681,
    17.95347, 17.90477, 18.29664, 18.37427, 17.97545, 20.12551, 21.45054,
    19.43811, 18.42702,
  17.87595, 17.88132, 17.78368, 17.99218, 17.8455, 17.73461, 17.75932,
    17.77588, 17.84851, 17.99802, 18.6474, 19.09389, 19.07485, 18.58008,
    18.44008, 18.40498, 17.93438, 17.89975, 18.24315, 18.82594, 18.8513,
    18.10386, 17.88547, 18.45581, 21.44535, 21.70263, 22.05844, 25.54354,
    21.14854, 19.32026,
  17.96774, 17.96612, 17.89516, 18.01465, 17.88813, 17.76886, 17.76608,
    17.82857, 17.94361, 18.07029, 18.16815, 18.65208, 19.12614, 19.35115,
    19.23191, 18.4604, 18.23116, 18.5206, 18.65516, 18.76477, 19.0206,
    19.73302, 20.47153, 19.77437, 24.79051, 28.0075, 24.56769, 25.67922,
    21.00467, 19.86893,
  17.83201, 17.84685, 18.01099, 18.08542, 18.2542, 18.61207, 18.62241,
    18.40429, 18.43078, 18.60896, 18.7292, 19.2308, 19.03381, 18.87266,
    19.60258, 20.10842, 19.54333, 18.65515, 18.4443, 18.21833, 20.40137,
    22.02633, 21.25635, 24.99223, 27.23743, 26.5962, 28.26244, 24.87073,
    20.63288, 19.1229,
  18.20173, 17.94686, 18.10325, 18.39643, 18.71367, 19.08273, 19.06287,
    18.72551, 19.20813, 19.80959, 19.90012, 19.55396, 18.98409, 19.01028,
    19.85315, 20.55572, 19.16872, 17.92714, 18.05352, 21.98635, 24.03633,
    20.75064, 20.36075, 23.42388, 25.10828, 24.53582, 24.73156, 24.55141,
    24.1983, 20.06909,
  18.21134, 18.03619, 18.61759, 19.55786, 19.7307, 19.33961, 19.29211,
    19.13721, 19.08639, 19.26675, 18.93668, 20.04819, 21.62504, 21.84698,
    21.13513, 25.2488, 29.72131, 24.47816, 20.72398, 24.27906, 23.13794,
    19.25193, 20.02621, 20.86472, 23.73469, 23.35485, 23.9495, 34.31649,
    32.93882, 20.03094,
  18.05056, 18.26937, 19.19271, 20.30802, 20.52898, 19.81736, 20.18161,
    21.61367, 21.60808, 21.43493, 21.95846, 22.1442, 21.83712, 21.50634,
    25.126, 32.10891, 31.77504, 24.47083, 21.87748, 22.09254, 20.44232,
    19.39248, 20.00419, 22.32603, 24.09499, 21.4215, 28.96689, 44.75159,
    35.71494, 18.603,
  18.20943, 18.5392, 19.56121, 20.54362, 20.26675, 21.49175, 23.68341,
    22.7991, 21.67639, 21.82468, 22.23713, 21.08274, 19.54334, 19.30204,
    22.85859, 25.9876, 23.9233, 21.56162, 20.51226, 20.32202, 19.81936,
    19.5339, 20.56304, 23.29953, 23.28837, 20.70294, 34.99226, 43.03128,
    26.35379, 18.55637,
  19.3466, 19.56889, 20.69246, 20.70494, 20.85056, 23.64055, 23.68023,
    21.40263, 21.29391, 21.57495, 20.91338, 19.5965, 18.76341, 22.26227,
    24.46758, 21.80278, 21.90428, 23.32848, 23.04884, 21.09817, 19.40707,
    20.42967, 24.46173, 25.60273, 22.53186, 22.3787, 31.86151, 31.36794,
    20.62069, 18.7326,
  21.42463, 22.05116, 24.28788, 26.1137, 26.28253, 23.78757, 20.47348,
    20.1698, 20.4608, 19.75349, 20.32284, 23.2107, 24.86538, 25.80308,
    25.44327, 24.57385, 24.9467, 25.80642, 25.2349, 23.71292, 22.98085,
    24.13017, 26.28072, 25.07758, 27.87911, 36.07572, 32.54271, 23.05768,
    19.65689, 18.06617,
  26.83447, 31.77994, 31.31736, 26.78817, 26.99707, 25.5701, 22.33152,
    23.91518, 24.89529, 30.15, 33.45016, 26.4914, 24.42397, 23.77371,
    22.74065, 24.01382, 25.64864, 25.74701, 24.39894, 24.15229, 26.73356,
    27.05718, 24.05908, 21.76889, 26.76773, 33.0306, 27.10193, 19.5341,
    18.40608, 17.78917,
  41.63475, 35.1496, 31.88261, 30.77761, 29.93162, 26.79744, 30.22737,
    30.18739, 26.71925, 32.15357, 33.05027, 22.38491, 22.45072, 23.72505,
    23.08115, 23.6496, 23.36757, 23.28277, 22.63399, 23.2805, 27.13118,
    26.16006, 21.50071, 24.20741, 26.9009, 22.26697, 18.79465, 18.60689,
    18.48652, 17.94135,
  52.87446, 40.75658, 43.6707, 49.8396, 51.71865, 49.93356, 42.2448,
    29.63622, 29.23984, 28.82119, 25.49014, 20.20359, 24.96643, 27.03063,
    24.50152, 23.75973, 23.65936, 22.76953, 22.22924, 25.26517, 27.87213,
    24.36687, 21.17021, 27.4869, 29.52138, 20.88363, 18.4289, 18.84077,
    19.04413, 18.25087,
  60.68673, 59.40761, 61.86897, 65.67478, 66.13268, 61.16505, 48.50943,
    43.5895, 36.56631, 30.61998, 35.60218, 36.45183, 39.80606, 40.59912,
    36.62656, 29.09969, 24.30951, 25.74781, 27.67471, 29.49418, 26.88457,
    25.35975, 27.66321, 26.14752, 23.19234, 19.48088, 18.53979, 18.48723,
    18.98345, 18.31544,
  43.52494, 45.73377, 50.96887, 57.83813, 59.49047, 52.90687, 53.18661,
    54.76588, 42.38796, 42.50264, 45.82645, 38.93666, 33.74969, 38.86694,
    39.83102, 29.04637, 27.83426, 28.09319, 30.67882, 31.94721, 28.81383,
    27.15363, 25.80365, 21.76995, 19.002, 19.39431, 18.69479, 18.28911,
    18.40472, 18.04645,
  28.96503, 32.84173, 38.02999, 40.79066, 38.32465, 36.41146, 39.60432,
    36.95395, 33.88958, 36.49979, 36.17009, 29.54733, 25.94236, 31.28333,
    30.85522, 28.05742, 29.89058, 27.83027, 28.29635, 29.00361, 25.79729,
    23.23601, 20.11843, 19.38036, 19.46926, 19.27605, 18.86532, 18.47621,
    18.26113, 17.92311,
  26.83485, 28.05615, 28.0725, 26.09323, 24.19592, 24.9582, 26.42918,
    25.94352, 26.92833, 27.88088, 25.04972, 25.62386, 28.91108, 27.80497,
    27.80066, 28.42588, 28.77082, 26.23145, 26.98643, 26.67132, 21.17577,
    20.64546, 19.85574, 19.39484, 19.23891, 19.26532, 18.80768, 18.28144,
    18.18335, 17.91532,
  23.23808, 22.60192, 20.99065, 20.31128, 20.70114, 22.01999, 22.90653,
    23.73676, 24.29608, 22.8871, 22.69858, 27.77115, 30.17118, 29.04607,
    32.34618, 31.13068, 27.07692, 24.01258, 26.88189, 25.79202, 20.40273,
    20.44305, 20.12785, 19.637, 18.89906, 19.00347, 18.63977, 18.00526,
    17.96641, 17.83175,
  21.90352, 21.11184, 19.25296, 18.9636, 19.47154, 20.01484, 20.57126,
    20.83424, 20.40926, 20.06924, 24.11141, 27.33021, 25.64815, 27.27579,
    29.65156, 28.69613, 27.04767, 26.02563, 28.56216, 26.59226, 22.1726,
    20.92274, 20.22413, 19.7773, 18.77892, 18.61442, 18.43771, 17.9795,
    17.89378, 17.79051,
  21.8795, 21.13279, 19.26201, 18.06532, 18.40331, 18.52159, 18.63152,
    18.65307, 18.59666, 21.57063, 25.31109, 24.3326, 23.08061, 24.14288,
    24.57553, 24.25956, 25.43424, 27.00922, 27.87005, 27.72891, 25.44904,
    22.62394, 20.4307, 19.86088, 19.10531, 18.57176, 18.34204, 18.01309,
    17.87732, 17.79175,
  21.02864, 20.77535, 19.16283, 17.89676, 17.88945, 17.96003, 17.8178,
    17.77979, 19.00596, 23.32378, 24.41861, 21.98478, 23.04824, 23.49818,
    22.90237, 22.30589, 22.69734, 23.40025, 24.07215, 24.72684, 25.30484,
    24.22071, 21.6783, 20.47883, 19.55389, 18.80858, 18.32291, 18.00182,
    17.89184, 17.79829,
  21.29465, 20.38449, 19.04924, 18.26612, 18.00891, 17.53681, 17.56818,
    18.06067, 20.49258, 23.52155, 22.41678, 20.78894, 22.26921, 22.6003,
    22.03951, 21.56811, 21.19813, 21.16717, 21.85505, 22.00025, 23.10996,
    23.23049, 22.28803, 22.35991, 20.95404, 19.1771, 18.3205, 18.04836,
    17.90779, 17.80204,
  21.49748, 20.53612, 18.92146, 18.16661, 18.5628, 18.77639, 18.94634,
    19.00342, 21.3293, 22.60435, 20.65289, 20.3287, 21.37875, 21.57409,
    21.13194, 21.32752, 21.27411, 20.70786, 20.62915, 20.58083, 21.66989,
    21.44494, 20.67852, 22.49817, 22.49208, 19.91464, 18.50317, 18.47395,
    18.16201, 17.82888,
  21.24546, 20.54239, 19.40994, 19.10015, 19.64134, 20.3306, 21.51802,
    22.39106, 23.48946, 21.71113, 19.64493, 20.49102, 21.50616, 21.98358,
    21.66726, 21.88427, 22.2676, 21.39866, 20.34821, 20.40184, 20.8203,
    20.38478, 19.80168, 20.54036, 21.75804, 21.43093, 19.83688, 18.93751,
    18.55713, 17.93186,
  21.27558, 20.99582, 19.53272, 19.41955, 20.58004, 21.60905, 22.20401,
    22.89398, 24.30755, 21.92077, 19.43114, 20.71553, 21.83985, 22.48231,
    22.55168, 22.59517, 22.48564, 22.02913, 21.03832, 20.46609, 20.33565,
    20.12381, 20.08134, 19.65455, 19.85038, 21.46801, 21.27606, 19.75154,
    19.52761, 18.37497,
  21.44058, 22.35152, 21.53457, 20.96642, 21.33844, 21.60225, 22.4023,
    23.51418, 22.99851, 21.08586, 19.70687, 21.04811, 22.37689, 22.59923,
    22.28158, 22.27581, 21.84692, 21.72109, 21.4238, 20.64795, 20.59905,
    20.62199, 19.84596, 19.26833, 19.26519, 20.23721, 21.67493, 20.56766,
    19.65796, 18.3875,
  22.55532, 23.72792, 22.9106, 21.94053, 21.22733, 20.61024, 22.86836,
    24.05094, 21.12794, 19.48685, 20.19386, 21.66916, 22.71603, 22.47158,
    21.84968, 21.61195, 21.26098, 21.31613, 21.17776, 20.55673, 20.72536,
    21.56161, 21.31878, 20.68398, 20.76118, 21.08171, 23.31171, 22.51356,
    19.33118, 17.82571,
  24.20467, 24.65665, 21.98369, 21.51625, 21.7335, 21.50331, 22.79462,
    21.94429, 18.79177, 18.7578, 20.29617, 21.69527, 22.26589, 22.12729,
    22.106, 21.68725, 20.95886, 20.85403, 21.35391, 21.70712, 22.08612,
    22.33193, 22.00486, 21.45895, 21.7173, 21.85821, 22.85178, 24.5753,
    22.03638, 18.38868,
  23.02464, 21.62139, 21.33007, 22.93796, 23.59898, 23.70799, 22.97921,
    19.76811, 17.886, 18.83881, 19.65143, 20.38258, 20.8588, 21.23059,
    21.86613, 21.97373, 21.74315, 22.03404, 22.09525, 21.95976, 22.0141,
    21.49648, 20.54622, 20.11625, 20.56415, 21.05206, 21.20603, 21.89388,
    22.35994, 19.18302,
  21.74829, 20.98507, 21.72181, 22.53453, 23.03289, 24.38611, 23.781,
    19.76913, 17.92694, 19.2043, 20.31878, 21.36226, 22.17422, 22.45791,
    22.59079, 22.74908, 22.15918, 21.66655, 21.33547, 20.48724, 19.96701,
    19.83605, 19.45743, 19.2867, 19.4831, 20.17579, 20.36492, 19.64262,
    19.45612, 18.27814,
  18.55335, 18.60394, 18.6154, 18.61182, 18.59816, 18.59865, 18.61012,
    18.63352, 18.66829, 18.69674, 19.46405, 19.62794, 18.72508, 18.91301,
    19.10559, 18.80124, 18.71723, 18.72461, 18.69681, 19.17201, 19.49313,
    19.07327, 19.02905, 19.44855, 19.47129, 19.05328, 21.36118, 23.42415,
    20.86681, 19.67877,
  18.81073, 18.89108, 18.70889, 18.96713, 18.80025, 18.63111, 18.67156,
    18.70601, 18.7672, 18.97685, 19.66983, 20.2227, 20.27076, 19.75073,
    19.51487, 19.52502, 18.89569, 18.86048, 19.32917, 20.0483, 20.045,
    19.19012, 18.92953, 19.68803, 22.94423, 24.23809, 23.98454, 28.75691,
    22.94686, 20.73717,
  18.90453, 18.93207, 18.82681, 18.97006, 18.83339, 18.66745, 18.66347,
    18.75972, 18.89694, 19.04824, 19.21877, 19.76199, 20.29548, 20.59735,
    20.53596, 19.58472, 19.25572, 19.67577, 19.81864, 19.96795, 20.27603,
    21.23297, 22.12965, 21.57439, 26.94925, 32.25657, 27.91963, 29.58423,
    22.96717, 21.44097,
  18.77483, 18.77682, 18.94221, 19.08064, 19.32198, 19.75866, 19.72182,
    19.42505, 19.4529, 19.69197, 19.88815, 20.46922, 20.32614, 19.98538,
    20.92887, 21.60015, 21.02759, 19.86233, 19.51658, 19.29937, 21.82565,
    24.04099, 23.05135, 27.70194, 31.00524, 29.90671, 33.31524, 28.44083,
    22.60723, 20.57201,
  19.19752, 18.87402, 19.09708, 19.4511, 19.87776, 20.24675, 20.1457,
    19.80123, 20.39948, 21.35901, 21.63913, 21.04779, 20.14572, 20.31213,
    21.34079, 21.96966, 20.45688, 18.85589, 19.07595, 23.84945, 26.96025,
    22.39106, 22.03535, 25.52522, 27.84929, 27.30677, 27.92922, 28.37253,
    27.95011, 21.94323,
  19.16527, 18.97405, 19.69732, 20.82419, 21.16348, 20.69363, 20.41479,
    20.25391, 20.23794, 20.60241, 20.3659, 21.5655, 23.63138, 23.82211,
    23.06352, 27.70309, 33.82673, 27.54303, 22.57763, 26.63973, 25.6002,
    20.58355, 21.49663, 22.67601, 25.8344, 25.85758, 26.22773, 39.41951,
    39.0079, 21.79499,
  19.00794, 19.29382, 20.37198, 21.67126, 22.1359, 21.39549, 21.43858,
    23.33521, 23.69049, 23.58881, 24.19466, 24.38066, 23.78107, 23.29341,
    27.37877, 36.05738, 35.90271, 26.88355, 23.84629, 24.20443, 22.10634,
    20.68966, 21.4745, 24.26087, 26.44658, 23.74781, 31.04824, 49.84309,
    41.95466, 20.003,
  19.15733, 19.6093, 20.82463, 22.00595, 21.77833, 23.18207, 25.8967,
    25.01105, 23.64151, 24.01103, 24.38936, 23.00121, 20.90148, 20.71605,
    24.80993, 28.8391, 26.16799, 23.44418, 22.13239, 21.93177, 21.28764,
    20.87913, 22.23755, 25.51986, 25.59141, 22.95363, 37.61882, 49.03807,
    29.60166, 19.80833,
  20.56646, 20.81722, 21.95886, 22.07885, 22.42429, 26.1589, 26.43386,
    23.24124, 23.1759, 23.65012, 22.83566, 21.01519, 19.93028, 23.94098,
    27.46822, 24.15786, 23.4979, 25.47243, 25.31321, 23.0231, 20.76412,
    22.17056, 27.01958, 28.58914, 24.47628, 24.67464, 34.87439, 35.77575,
    22.3101, 19.90979,
  23.01328, 23.57367, 26.20732, 29.18324, 29.21011, 26.54234, 22.2368,
    21.65347, 21.86775, 21.20267, 21.70547, 25.11522, 27.01802, 28.17808,
    27.81359, 26.81536, 27.30215, 28.33719, 27.71105, 25.75555, 25.13146,
    26.55931, 28.89464, 27.62087, 30.61895, 40.90827, 37.65292, 25.17072,
    20.8654, 19.07406,
  30.27915, 35.80665, 36.76007, 30.34043, 30.13215, 28.78164, 25.49936,
    26.87498, 28.02576, 32.12805, 36.9033, 29.20949, 26.61579, 25.87356,
    24.9646, 26.43917, 28.46922, 28.67459, 27.09485, 26.18314, 29.25172,
    29.74256, 26.17724, 23.42952, 29.0181, 36.34687, 30.06668, 20.69977,
    19.46782, 18.69661,
  47.19722, 39.8623, 36.65258, 33.76539, 33.64661, 28.63383, 32.77643,
    33.49811, 29.79392, 35.0094, 35.92973, 23.90263, 24.14648, 25.88629,
    25.24888, 26.28835, 25.92812, 25.95342, 25.0394, 25.50664, 29.80886,
    28.68848, 22.99495, 25.83239, 29.79957, 24.60847, 20.01455, 19.63,
    19.50433, 18.89772,
  61.82767, 48.08172, 49.54914, 55.861, 57.89722, 55.5205, 49.29382,
    42.70905, 49.53279, 37.04139, 28.32276, 24.30176, 29.00231, 29.47568,
    27.52959, 26.29409, 26.25388, 25.2473, 24.26425, 27.83333, 31.0612,
    26.2243, 22.54066, 29.26692, 32.79591, 22.60173, 19.40374, 19.8904,
    20.11436, 19.28862,
  69.8915, 59.84964, 62.3381, 69.02055, 73.23997, 73.09835, 63.97295,
    63.11485, 53.93156, 37.96564, 39.54891, 39.16839, 41.85331, 44.77389,
    41.74664, 31.92352, 27.19704, 28.98647, 31.53821, 33.93791, 30.4081,
    26.73329, 30.02671, 28.70007, 25.22726, 20.66479, 19.54425, 19.5174,
    20.01493, 19.39876,
  59.16079, 70.18026, 75.11594, 82.42209, 82.64853, 71.20369, 67.71246,
    70.17921, 49.02476, 47.98559, 56.21027, 55.92878, 58.71474, 54.22028,
    43.58031, 33.72969, 31.75373, 32.25087, 35.38437, 36.83873, 31.72848,
    29.54805, 28.41356, 24.0013, 20.21818, 20.46252, 19.71677, 19.30195,
    19.38177, 19.06245,
  45.66332, 56.37728, 62.48938, 62.80214, 53.1976, 54.84578, 62.67677,
    45.33127, 48.92635, 57.67258, 50.35262, 43.11754, 42.84399, 41.54543,
    34.21861, 32.46487, 34.41219, 31.96953, 31.586, 32.63675, 28.23726,
    25.48377, 22.23924, 20.93479, 20.71252, 20.38158, 19.86357, 19.49015,
    19.224, 18.8875,
  36.27443, 38.44815, 39.42684, 35.61221, 31.27419, 36.88528, 41.72285,
    35.24921, 40.77316, 44.02992, 34.08775, 30.7219, 34.12173, 31.36959,
    31.72226, 32.31187, 33.14753, 29.85581, 29.7698, 30.64713, 23.31771,
    22.24858, 21.32728, 20.87562, 20.49164, 20.29924, 19.83506, 19.3143,
    19.16788, 18.90049,
  29.80065, 30.19153, 27.72105, 25.98603, 26.529, 28.32889, 29.51514,
    31.00275, 30.55807, 28.24076, 27.10766, 32.19275, 34.97055, 32.45908,
    37.42417, 36.12969, 31.07486, 26.64204, 29.85386, 29.47712, 21.98619,
    21.98698, 21.57584, 21.06933, 20.04964, 19.98874, 19.68052, 19.00726,
    18.95143, 18.81282,
  28.21071, 27.45385, 24.43883, 23.69108, 24.38128, 25.13517, 25.89476,
    25.87007, 24.99318, 23.67351, 27.56143, 31.49038, 28.8592, 30.48648,
    34.41108, 33.08997, 30.68407, 28.69604, 31.955, 29.82614, 23.95945,
    22.54026, 21.7417, 21.14673, 19.85889, 19.59616, 19.44711, 18.95918,
    18.84505, 18.73534,
  27.6755, 26.46102, 23.95725, 22.46585, 22.97365, 23.20139, 23.3384,
    23.24474, 22.62926, 25.23147, 29.14798, 27.2909, 25.14038, 26.75639,
    27.89426, 27.69361, 28.84701, 30.52804, 31.2075, 30.80163, 27.65983,
    24.57974, 22.0313, 21.17682, 20.17501, 19.55856, 19.33255, 19.00932,
    18.83044, 18.73589,
  26.17633, 25.74539, 23.67575, 22.08845, 22.1257, 22.30893, 22.18471,
    21.8601, 22.71436, 27.08204, 27.99944, 24.06579, 25.13047, 25.8908,
    25.38977, 24.90236, 25.56487, 26.50795, 26.78259, 27.41971, 28.01372,
    26.97092, 23.413, 21.87163, 20.69699, 19.90965, 19.35962, 19.02335,
    18.84796, 18.74575,
  26.47834, 25.17113, 23.45669, 22.44038, 22.29285, 21.70712, 21.64675,
    21.8998, 24.3754, 27.47687, 25.48386, 22.69636, 24.42052, 24.88523,
    24.30283, 23.75945, 23.45868, 23.32931, 24.11453, 24.39476, 25.71985,
    26.05191, 23.93358, 24.13082, 22.52766, 20.48198, 19.39882, 19.07643,
    18.85571, 18.75164,
  26.60024, 25.18515, 23.2824, 22.31856, 22.89212, 23.0201, 23.06489,
    22.84804, 25.33634, 26.58852, 23.32993, 22.36366, 23.50023, 23.68882,
    23.20755, 23.45767, 23.4052, 22.71449, 22.64197, 22.58995, 23.82185,
    23.74862, 22.18097, 24.33564, 24.40582, 21.44497, 19.58054, 19.55904,
    19.14639, 18.78071,
  26.20928, 25.11966, 23.94777, 23.53244, 24.0764, 24.53834, 26.02291,
    27.37989, 28.55676, 25.78197, 22.23797, 22.70283, 23.64196, 24.20907,
    23.85736, 24.06385, 24.52132, 23.56607, 22.27575, 22.30614, 22.90844,
    22.21285, 21.18747, 22.20082, 23.59563, 23.20736, 21.29253, 20.09542,
    19.60861, 18.92225,
  26.11939, 26.26356, 24.15217, 23.55066, 24.93151, 26.34757, 27.30631,
    28.30608, 29.63802, 26.2856, 22.07168, 23.04889, 24.08578, 24.905,
    24.97864, 25.07602, 24.93851, 24.30102, 22.9819, 22.26148, 22.09963,
    21.63498, 21.62743, 21.27332, 21.33187, 23.06701, 22.86939, 21.03582,
    20.6916, 19.53948,
  26.56153, 28.27205, 26.74905, 25.62761, 26.14527, 26.78481, 27.99515,
    29.40326, 28.19095, 25.38357, 22.49745, 23.4611, 24.78719, 25.13825,
    24.76306, 24.85099, 24.30674, 23.89961, 23.30994, 22.20659, 22.14887,
    22.25935, 21.4356, 20.60718, 20.43805, 21.55831, 23.16961, 22.07057,
    20.84973, 19.60559,
  27.93346, 29.85941, 28.45014, 26.88859, 26.36323, 25.83797, 28.97317,
    30.64307, 26.21535, 23.31527, 23.10756, 24.20727, 25.13057, 24.9117,
    24.26849, 24.01719, 23.51079, 23.31254, 22.97989, 22.06758, 22.36912,
    23.35984, 22.99406, 22.03059, 22.00789, 22.49387, 24.90521, 24.29232,
    20.61627, 18.89969,
  29.89892, 31.24815, 27.1885, 26.18484, 26.85164, 26.91618, 28.96143,
    28.23881, 23.43023, 22.27322, 23.14832, 24.15477, 24.58904, 24.4554,
    24.51187, 24.06059, 23.02427, 22.69503, 23.08783, 23.44048, 24.16325,
    24.61479, 23.99676, 23.10136, 23.15132, 23.53978, 24.69898, 26.46615,
    23.77623, 19.57024,
  28.68509, 26.95575, 26.52501, 30.02033, 30.50169, 29.7697, 29.51723,
    25.53707, 22.18926, 22.33013, 22.38151, 22.56743, 22.88682, 23.36423,
    24.24803, 24.34866, 23.78249, 23.99895, 24.14374, 23.9852, 24.20994,
    23.62757, 22.27986, 21.57397, 22.01922, 22.71162, 23.01029, 23.72195,
    24.03834, 20.60779,
  26.89199, 25.84306, 27.78004, 30.7987, 30.77879, 31.12061, 30.3181,
    25.09777, 21.91636, 22.56635, 22.79364, 23.29244, 24.03799, 24.49181,
    24.85712, 25.03452, 24.27717, 23.66563, 23.26047, 22.24165, 21.59689,
    21.30087, 20.78111, 20.54444, 20.8342, 21.6535, 21.99417, 21.16494,
    20.72804, 19.44137,
  26.05893, 26.13781, 26.17008, 26.19554, 26.17863, 26.17808, 26.18541,
    26.2681, 26.40429, 26.6724, 28.17033, 28.70354, 26.65204, 26.78035,
    26.95163, 26.45913, 26.32408, 26.39818, 26.51688, 27.2901, 27.98936,
    27.4771, 27.76965, 28.9732, 29.93301, 30.3727, 34.45018, 38.08757,
    31.01693, 28.06317,
  26.71883, 26.99651, 26.48628, 27.05274, 26.73756, 26.34464, 26.45936,
    26.5666, 26.81843, 27.3155, 28.29569, 29.39028, 29.90873, 28.79728,
    27.75084, 28.05087, 26.8636, 27.00833, 28.09097, 29.24145, 28.7572,
    27.57937, 28.43033, 31.99216, 38.84449, 41.65854, 38.59347, 44.99107,
    33.59705, 29.70364,
  26.79894, 26.8799, 26.7006, 26.83989, 26.62063, 26.44745, 26.49073,
    26.6932, 26.93506, 27.1827, 27.59913, 28.53493, 29.38112, 30.02464,
    30.05682, 28.22589, 27.91339, 28.88507, 28.99867, 29.44181, 31.08304,
    33.54062, 36.08804, 40.08185, 47.56376, 53.11432, 46.24797, 46.12207,
    33.89021, 31.20458,
  26.6673, 26.71597, 27.0403, 27.48775, 28.02408, 28.95495, 28.88668,
    28.13228, 28.26048, 28.95241, 29.5048, 30.18228, 29.85647, 29.04762,
    30.9163, 32.37151, 31.388, 29.03872, 29.05003, 30.55713, 36.49952,
    41.0157, 39.81705, 48.04897, 54.83415, 50.09341, 54.57886, 44.0891,
    33.64227, 29.49285,
  27.61097, 26.95055, 27.58287, 28.37761, 29.33805, 29.7378, 29.34621,
    29.02708, 30.43677, 31.98716, 31.48567, 30.34552, 29.47775, 30.16506,
    31.65993, 32.18841, 30.38103, 28.5929, 31.36772, 39.90059, 45.38213,
    37.69781, 37.68457, 41.56494, 45.39643, 44.62389, 42.91402, 46.1213,
    43.3073, 30.88185,
  27.38356, 27.55013, 29.16632, 31.39518, 31.54453, 30.33182, 30.39478,
    30.05527, 29.4633, 29.83082, 29.87661, 32.93279, 38.04701, 37.04226,
    38.82795, 47.27926, 51.98265, 46.63252, 40.05645, 44.53738, 41.59243,
    33.80799, 35.76787, 38.5149, 41.78848, 42.05565, 45.45407, 63.51577,
    58.48311, 30.22682,
  27.5544, 28.78944, 30.94505, 33.26684, 33.09122, 31.62548, 33.27318,
    37.14134, 38.21146, 38.06318, 39.72464, 39.80356, 37.64277, 38.37396,
    45.65815, 56.31822, 53.77291, 45.19208, 39.43721, 39.15449, 35.60822,
    33.30053, 35.2853, 40.73906, 44.93582, 44.52569, 53.98541, 70.22404,
    58.75761, 28.20567,
  28.0797, 29.84741, 32.26132, 34.27967, 33.67321, 37.56688, 44.14405,
    40.21926, 36.67237, 37.65428, 37.52777, 35.33614, 32.85666, 34.59706,
    39.64215, 44.67292, 42.59607, 39.70815, 34.76862, 34.27363, 33.0315,
    32.84225, 36.42826, 42.52686, 44.39737, 44.62663, 59.42557, 67.61478,
    44.91071, 28.33633,
  30.2331, 30.82891, 33.96946, 35.52351, 36.03756, 41.14425, 40.41955,
    35.78706, 36.19484, 36.55906, 34.6843, 31.81676, 31.80251, 40.50938,
    48.00418, 40.99814, 38.38616, 41.16887, 41.40575, 37.26617, 33.15727,
    37.18612, 45.56631, 48.84832, 42.1778, 46.76678, 59.45758, 55.2448,
    34.56236, 28.23978,
  35.39997, 42.45227, 44.6235, 45.55913, 45.72587, 42.04702, 31.73703,
    31.29636, 30.49455, 30.39522, 31.88577, 40.06741, 47.35945, 47.30527,
    43.63215, 42.93587, 44.18826, 46.37002, 44.50543, 38.90378, 39.85406,
    42.1117, 44.94683, 46.33364, 55.43633, 68.97791, 60.07218, 36.66443,
    29.30355, 26.67723,
  48.17756, 54.50926, 54.43701, 48.14637, 47.96547, 43.29333, 35.26011,
    39.30774, 44.84681, 51.83603, 56.86887, 43.89351, 40.02384, 38.83213,
    37.7488, 40.51675, 43.25423, 43.38723, 41.09288, 38.72167, 43.09149,
    44.01151, 39.39811, 37.76154, 45.27277, 50.43164, 39.5418, 28.01473,
    27.36799, 26.21192,
  67.03532, 53.23388, 51.68742, 51.82489, 50.72411, 42.63752, 50.02808,
    53.06511, 49.05221, 51.03097, 47.31733, 34.19344, 35.372, 37.82167,
    38.41164, 40.59366, 40.02736, 39.35082, 38.12682, 39.68927, 43.59303,
    41.44687, 34.06338, 38.97383, 44.68219, 34.80527, 27.60427, 27.72005,
    27.46706, 26.55125,
  78.66409, 64.92806, 76.48052, 85.32336, 87.19743, 81.1573, 68.69037,
    52.97778, 54.24915, 43.88441, 36.16825, 32.04935, 39.60619, 44.63132,
    43.51947, 40.95779, 40.58762, 38.71612, 38.2847, 45.09133, 45.99775,
    37.79788, 33.96312, 40.92192, 45.77874, 31.17793, 27.33282, 28.18272,
    28.35941, 27.21001,
  86.21973, 100.3378, 104.3541, 107.4313, 100.1475, 91.00391, 78.7775,
    72.65337, 58.1218, 47.70879, 58.08147, 60.02925, 65.96216, 67.83384,
    62.41778, 50.33675, 42.42166, 45.21105, 49.31572, 51.71409, 44.74539,
    38.27348, 43.85632, 39.14991, 33.65149, 28.99239, 27.66162, 27.53097,
    28.05578, 27.30888,
  86.73272, 89.04594, 91.67935, 87.8623, 76.69916, 73.44357, 85.29932,
    81.27993, 67.4398, 73.12427, 76.43623, 67.0888, 61.539, 67.32858,
    66.11681, 52.92536, 51.03376, 53.30661, 57.97473, 58.56961, 48.01236,
    44.75154, 40.59552, 32.35336, 28.42661, 28.78277, 27.82615, 27.24265,
    27.19662, 26.76544,
  83.16208, 83.3884, 78.63875, 69.72927, 64.62576, 67.64789, 76.59082,
    77.72304, 75.10373, 64.42883, 64.92605, 54.7836, 49.15411, 56.0761,
    54.50547, 52.43518, 56.11703, 54.86865, 56.51205, 54.21154, 41.31396,
    36.56103, 32.00692, 29.54477, 29.156, 28.63429, 27.89907, 27.43146,
    27.02386, 26.55636,
  72.80794, 66.11781, 57.5627, 53.58216, 53.92882, 55.33319, 60.29668,
    65.3604, 59.31734, 55.06079, 47.11697, 46.05128, 53.48203, 53.95691,
    51.66935, 53.29493, 53.54626, 49.41873, 50.40241, 49.13459, 33.33708,
    30.78353, 30.10534, 29.87663, 28.92792, 28.56957, 27.91447, 27.07385,
    26.87127, 26.55064,
  54.03172, 48.22083, 42.74478, 43.33623, 45.85255, 50.02411, 52.10793,
    51.12488, 48.06903, 43.74851, 42.70666, 52.71644, 56.43991, 57.28294,
    60.48721, 56.94165, 48.84181, 44.29556, 49.43468, 45.46444, 30.96455,
    31.73404, 31.24889, 30.1675, 28.20331, 28.10496, 27.76762, 26.66429,
    26.55607, 26.37318,
  45.13841, 42.43324, 37.86211, 37.41762, 41.3474, 44.51908, 43.4338,
    40.63672, 37.30264, 35.94183, 44.53151, 52.16006, 48.54283, 52.73609,
    54.36249, 48.87365, 47.63671, 50.62103, 53.60056, 47.07956, 35.95966,
    34.23572, 32.13085, 30.23065, 27.91453, 27.5928, 27.34154, 26.57759,
    26.43275, 26.3013,
  42.03634, 41.17199, 36.54835, 35.01785, 37.9247, 38.02678, 35.41756,
    32.79076, 32.10315, 39.98261, 48.81857, 45.39584, 43.2917, 45.52065,
    44.03141, 41.05218, 43.796, 50.05676, 51.99421, 50.13976, 43.91254,
    37.74134, 32.59606, 30.34155, 28.48996, 27.61302, 27.18023, 26.68448,
    26.39926, 26.30106,
  39.13891, 39.76167, 34.92143, 33.19917, 34.15522, 32.93495, 30.56711,
    29.94394, 34.18348, 44.40992, 46.47283, 38.76068, 40.72951, 40.50233,
    38.65648, 38.04426, 40.85662, 44.57684, 46.84725, 46.86359, 43.45494,
    39.74944, 34.93537, 31.42636, 29.25655, 28.23099, 27.2515, 26.75828,
    26.4502, 26.31387,
  39.82417, 37.82734, 33.84624, 32.42109, 31.84874, 29.40333, 29.22035,
    31.02611, 38.04517, 44.36486, 39.924, 34.80247, 37.01051, 36.19786,
    35.97931, 37.3167, 39.57296, 41.35798, 42.40515, 41.24483, 39.19735,
    38.01046, 36.11757, 35.50489, 32.55011, 29.24227, 27.3671, 26.9036,
    26.49563, 26.33284,
  39.55389, 38.02189, 32.73824, 30.49884, 31.22563, 31.89632, 32.91425,
    33.85098, 39.25923, 41.26602, 34.07969, 32.23582, 33.09809, 33.20877,
    34.29257, 37.44279, 39.84779, 39.34482, 38.20958, 36.46304, 35.84986,
    35.63493, 34.135, 36.07655, 35.60872, 30.94008, 27.65168, 27.71003,
    26.99604, 26.39215,
  38.80964, 36.99823, 34.2543, 32.95877, 33.97203, 35.7131, 38.21018,
    38.09786, 41.66624, 39.25257, 30.947, 31.11162, 32.31569, 34.42283,
    36.50256, 39.34751, 41.28314, 39.51191, 36.39829, 34.86243, 34.19286,
    33.50228, 32.98492, 33.83643, 34.78853, 33.63359, 30.53563, 28.45098,
    27.64111, 26.65281,
  37.13719, 38.88314, 33.45982, 31.81005, 34.29251, 36.54473, 37.67525,
    38.45186, 43.20719, 39.02696, 29.30821, 30.8436, 33.27597, 36.62844,
    39.17091, 41.28473, 41.35827, 39.50896, 35.98331, 33.26521, 33.28134,
    33.48998, 32.91888, 31.62034, 31.19676, 32.81092, 32.40625, 29.85115,
    29.05496, 27.62684,
  38.70183, 41.83821, 37.02748, 34.62416, 35.63717, 36.39267, 37.60337,
    40.871, 42.44622, 35.57271, 29.81685, 32.25759, 35.91749, 38.44546,
    39.36324, 40.55438, 39.83557, 37.85902, 35.02371, 32.49355, 33.85114,
    34.43172, 31.66923, 29.45191, 29.22201, 30.71721, 32.61703, 31.44271,
    29.27124, 27.71331,
  41.76889, 44.15559, 39.62442, 36.72511, 37.4971, 35.91102, 38.67807,
    41.48293, 38.60087, 31.40726, 31.51419, 34.79889, 37.6914, 38.47609,
    38.45735, 38.75594, 37.78549, 36.0811, 33.95401, 32.15606, 33.88697,
    35.45631, 33.79956, 31.6873, 31.39239, 32.27765, 35.25636, 34.69075,
    29.17498, 26.63361,
  44.82241, 45.9287, 38.71863, 37.72981, 39.92738, 38.60316, 40.82505,
    39.99049, 32.88052, 30.58647, 33.1669, 36.14164, 37.54815, 37.62322,
    38.32841, 38.1742, 36.24017, 34.63335, 33.87195, 34.31416, 36.82433,
    37.68776, 35.24263, 33.33101, 33.03216, 33.93975, 35.29186, 37.3867,
    33.96564, 27.79694,
  40.7641, 36.49095, 35.4126, 40.52814, 42.49012, 44.759, 43.78087, 36.84902,
    30.45297, 31.77117, 33.00722, 33.68809, 34.05616, 35.0152, 37.15261,
    38.00293, 37.21935, 36.7904, 35.6198, 34.89869, 36.18505, 35.18414,
    32.42473, 31.02399, 31.57433, 32.74584, 33.26572, 33.81312, 33.66504,
    29.36799,
  36.84164, 35.22585, 38.18416, 40.30983, 39.98882, 44.26067, 46.26552,
    36.60723, 31.14585, 33.31477, 34.14716, 34.87833, 35.8562, 37.13303,
    38.72807, 39.67132, 38.21622, 35.85095, 33.99265, 32.23351, 31.45807,
    30.54802, 29.68327, 29.35111, 29.89355, 31.03951, 31.46057, 30.43788,
    29.21184, 27.28508,
  28.3267, 28.57351, 28.85059, 29.16575, 29.25925, 29.53772, 29.98623,
    30.57508, 31.36424, 32.76223, 35.43516, 35.79845, 31.43237, 32.33614,
    32.62495, 31.08854, 31.34403, 32.53676, 34.20086, 37.20717, 39.18407,
    38.16023, 39.84819, 43.4455, 46.18531, 47.41498, 53.93118, 56.62828,
    37.13219, 31.39527,
  31.16874, 31.81601, 30.67641, 32.08911, 31.59684, 31.30442, 32.15627,
    32.97044, 34.01414, 35.33086, 37.2529, 39.60516, 40.62332, 37.81623,
    35.86252, 37.00786, 35.77816, 38.19827, 41.5631, 44.66046, 45.5724,
    46.22881, 49.49096, 56.78701, 63.71087, 61.02807, 55.58868, 59.69728,
    39.23607, 33.42841,
  29.68391, 29.87224, 30.11377, 30.60308, 30.8201, 31.2381, 31.76534,
    32.53755, 33.54301, 34.63938, 36.08432, 38.34602, 40.63669, 43.18671,
    44.94135, 43.41297, 46.1093, 50.53297, 53.91512, 59.41187, 67.61516,
    76.21853, 79.23352, 78.19191, 78.84719, 75.99864, 69.49087, 59.10714,
    40.06707, 35.69947,
  30.98688, 31.89184, 33.80084, 36.09233, 38.14388, 40.18082, 40.25707,
    39.73711, 41.03413, 42.97836, 44.23636, 45.82219, 46.98915, 48.26978,
    55.09367, 59.98321, 59.3342, 58.27799, 64.25824, 71.12299, 81.9328,
    86.00273, 79.08153, 84.56483, 85.55515, 82.72211, 76.98889, 56.44576,
    40.24625, 32.7803,
  35.86462, 35.50215, 38.39689, 40.63724, 42.32847, 41.99818, 41.46286,
    41.92832, 44.521, 46.76022, 46.47217, 47.86831, 50.38318, 54.93579,
    59.73917, 63.26788, 63.09805, 61.65065, 66.68442, 76.00002, 79.05281,
    67.70596, 68.77797, 75.78584, 82.3851, 83.10457, 73.89346, 78.01482,
    69.09076, 41.65531,
  36.76362, 39.35091, 43.28082, 47.26422, 46.27787, 43.79235, 45.00192,
    46.65814, 49.05643, 54.37037, 62.14164, 74.7692, 87.47958, 86.57936,
    88.62843, 93.55863, 97.52274, 89.64526, 78.00735, 77.48051, 69.57916,
    61.57744, 67.78923, 74.81501, 82.75269, 82.27014, 76.5352, 90.2106,
    78.98137, 39.26463,
  39.99091, 44.65374, 50.49131, 57.10148, 60.79392, 65.42116, 75.43484,
    86.55312, 90.01307, 90.62657, 91.6976, 86.3565, 76.88394, 77.34146,
    79.79284, 82.58844, 81.5003, 74.92818, 66.38921, 66.81677, 63.55926,
    63.42577, 69.61424, 78.44048, 79.97198, 70.24084, 72.07545, 82.42337,
    68.231, 31.23715,
  47.52548, 55.4571, 64.05, 73.1699, 78.11897, 87.71544, 95.10931, 80.84547,
    70.20217, 69.56532, 64.62164, 58.64721, 54.0293, 55.50771, 58.6286,
    63.59762, 66.47635, 65.49471, 58.34158, 59.44086, 59.56255, 62.97388,
    70.91394, 76.80153, 71.9866, 66.81992, 77.41208, 78.10093, 54.11129,
    32.03297,
  61.81043, 67.7132, 73.93893, 76.85934, 76.63014, 78.95295, 69.12083,
    62.77555, 63.76882, 63.46134, 61.56653, 60.38361, 64.54314, 78.74397,
    87.14998, 72.22911, 73.56644, 79.87681, 78.60526, 71.002, 69.05193,
    82.27626, 96.0191, 94.04576, 77.61622, 83.40884, 84.16855, 70.4149,
    40.06719, 31.58304,
  83.78056, 93.01974, 89.84365, 92.41484, 84.4436, 72.32765, 54.97116,
    62.65334, 66.19215, 76.043, 87.30267, 99.84254, 99.58191, 96.03902,
    91.54916, 97.91512, 102.1632, 99.91849, 92.27364, 89.14442, 97.28036,
    97.54898, 93.09413, 82.31167, 87.07206, 97.73647, 81.19939, 47.32554,
    31.76155, 28.10757,
  107.5721, 101.6215, 99.96021, 89.71909, 98.215, 98.96976, 96.8728,
    105.1228, 113.8129, 117.2079, 107.6572, 82.20551, 77.55763, 78.68419,
    81.81924, 88.3591, 92.16997, 90.63354, 86.82549, 86.32668, 96.90035,
    92.52032, 71.36183, 64.07993, 70.92989, 69.08278, 47.53043, 31.45987,
    30.15538, 27.8465,
  110.8028, 93.75023, 105.3943, 114.4494, 115.259, 102.1155, 105.7512,
    100.7617, 90.16117, 78.86459, 70.21602, 65.07322, 71.98683, 78.36665,
    80.7903, 81.28073, 78.91325, 77.04675, 73.73499, 74.95216, 83.63779,
    76.51783, 58.85854, 67.59301, 70.25758, 50.22216, 31.06946, 32.93615,
    31.04373, 28.85651,
  127.5563, 128.7589, 133.3056, 135.6388, 135.9315, 131.6396, 104.0184,
    91.38913, 94.71657, 72.37647, 70.99368, 73.92015, 85.82333, 94.46274,
    90.68676, 77.62242, 76.92424, 73.21198, 70.51882, 76.01279, 79.31129,
    68.42933, 60.37965, 59.68, 56.05339, 41.11103, 32.68328, 34.48788,
    33.26085, 30.41604,
  132.0901, 134.1599, 133.6574, 131.5591, 128.5247, 123.7305, 123.4838,
    123.8808, 106.9887, 110.8775, 123.6545, 119.6876, 126.05, 127.5887,
    113.3439, 93.06226, 90.66897, 94.62656, 98.54394, 92.26038, 77.08345,
    64.03729, 59.43773, 46.77971, 39.03699, 35.9838, 32.84377, 31.93328,
    31.7884, 30.24337,
  125.5386, 114.3093, 110.8172, 109.007, 110.306, 118.6011, 126.6444,
    127.6759, 125.4259, 126.4618, 126.1035, 124.026, 127.2641, 127.1573,
    121.3308, 117.3748, 106.5759, 104.2284, 103.1786, 91.09019, 63.5358,
    55.77081, 44.81145, 38.68198, 36.15641, 34.57841, 32.24914, 30.68971,
    29.73288, 28.81416,
  104.5445, 104.179, 107.3857, 110.5327, 115.1747, 125.3804, 128.806,
    127.4906, 121.8685, 120.265, 118.935, 110.8677, 106.5616, 118.1154,
    113.8255, 107.92, 104.1469, 91.63898, 83.28472, 69.85498, 47.33038,
    44.96274, 38.49828, 37.17627, 36.07313, 33.94661, 31.89948, 30.74381,
    29.50832, 28.59936,
  91.43961, 89.81931, 93.79226, 99.10285, 104.1918, 109.1012, 112.2225,
    112.847, 109.0613, 106.1608, 99.02217, 108.151, 121.4637, 112.5908,
    105.3435, 96.90913, 86.95603, 75.25096, 71.16849, 63.20488, 41.6689,
    42.88581, 39.02171, 37.14354, 35.55318, 34.29033, 31.71258, 29.60274,
    29.06517, 28.55764,
  75.69367, 80.33742, 81.59457, 86.23235, 89.45123, 93.04886, 94.65295,
    96.35599, 98.67159, 98.90278, 112.0714, 128.8192, 127.4676, 119.9151,
    112.3773, 93.23344, 72.86882, 64.77795, 69.66258, 61.59819, 43.1746,
    43.99456, 40.09961, 37.82717, 34.15703, 32.48119, 31.01882, 28.63964,
    28.40913, 28.1132,
  83.57709, 82.65894, 73.87389, 71.21785, 74.39519, 76.82051, 80.74387,
    86.50989, 91.27708, 100.3387, 114.7493, 114.1789, 95.39383, 93.94095,
    88.04459, 80.55167, 80.82652, 84.71611, 85.49576, 71.63008, 51.59863,
    45.2572, 40.3662, 36.86464, 32.66138, 31.0112, 30.0867, 28.54754,
    28.17727, 28.02846,
  82.0098, 76.47467, 65.97961, 60.22597, 64.35709, 69.06656, 75.57709,
    82.62465, 90.90958, 102.4437, 104.0497, 83.86452, 75.62931, 73.7303,
    71.11289, 71.70221, 77.28192, 84.04012, 82.57224, 75.48406, 61.3113,
    49.52947, 41.20916, 37.04885, 33.69983, 31.14633, 29.94121, 28.80337,
    28.14204, 28.02601,
  73.10365, 67.27463, 58.39098, 55.30328, 60.54002, 66.83747, 72.84451,
    78.41515, 84.13516, 88.73927, 80.00333, 64.51099, 69.43511, 69.97607,
    69.26712, 68.61742, 70.32338, 70.38219, 68.43784, 63.83369, 57.70896,
    54.08639, 46.6216, 40.31316, 36.08457, 32.68608, 29.96216, 28.79722,
    28.15858, 28.0575,
  70.64799, 61.8819, 57.11479, 56.93023, 61.89774, 63.83948, 68.7924,
    71.46419, 76.553, 77.49313, 66.22132, 59.5511, 66.18312, 67.07143,
    65.79632, 63.96364, 61.29728, 58.04599, 56.2909, 54.15104, 52.6909,
    51.26391, 49.47174, 48.26107, 42.0943, 34.26274, 30.07051, 29.13129,
    28.1912, 28.02094,
  65.85329, 61.3666, 56.54249, 57.46047, 65.52492, 69.55107, 70.02771,
    66.83133, 68.2492, 66.04345, 55.89558, 58.09306, 62.02547, 62.61143,
    59.86916, 58.51421, 56.27502, 51.13503, 49.02886, 48.51593, 48.05379,
    46.92691, 45.19379, 46.9229, 46.56229, 37.98486, 31.82026, 31.46478,
    29.46009, 28.13581,
  67.24298, 66.69107, 67.55263, 70.63062, 75.09593, 74.5255, 75.41258,
    72.62228, 72.85757, 64.43969, 55.35062, 61.29348, 64.15881, 64.88882,
    61.57483, 59.47692, 58.03902, 53.19624, 48.67797, 47.50384, 46.27338,
    44.37614, 42.99529, 43.23278, 44.8065, 44.08199, 38.32607, 32.98005,
    31.02672, 28.86978,
  71.29002, 74.18828, 70.1695, 70.91608, 73.77344, 72.30882, 70.18082,
    70.95897, 75.79745, 67.64886, 56.63284, 63.07077, 65.47427, 66.39006,
    64.09344, 62.55533, 58.7883, 54.83407, 50.60542, 46.47277, 45.72468,
    45.35146, 42.987, 41.04693, 41.01868, 43.79993, 43.4543, 37.9334,
    34.92554, 31.478,
  80.9397, 86.45285, 84.07561, 77.94016, 73.82979, 71.05939, 75.48937,
    80.61551, 76.32561, 65.61241, 62.07678, 66.31448, 68.54887, 66.96622,
    63.01644, 61.28946, 58.08304, 54.83838, 51.98779, 47.99835, 47.09868,
    45.57592, 41.47258, 39.39269, 40.25134, 42.59288, 44.87067, 41.31537,
    34.45035, 31.0146,
  91.66888, 93.41388, 82.07913, 75.27815, 72.1133, 70.30827, 79.02658,
    80.64183, 69.11753, 62.44246, 65.85104, 67.92086, 67.71515, 65.07697,
    61.89056, 59.31498, 55.76171, 52.90497, 50.43708, 47.63139, 48.78424,
    51.17033, 50.39003, 47.70337, 47.36627, 48.74323, 51.68727, 47.80627,
    34.6892, 28.86559,
  94.1647, 88.1211, 78.40707, 78.13439, 79.75735, 79.70534, 82.52577,
    75.43787, 63.20668, 64.35581, 66.73779, 67.23513, 66.38266, 63.94994,
    61.9716, 58.413, 53.98341, 52.79876, 54.918, 57.70135, 59.29423,
    57.79051, 53.70479, 51.67427, 51.29945, 52.3768, 53.04147, 54.30356,
    46.69376, 32.26225,
  80.31343, 76.15266, 81.67562, 89.3245, 92.205, 93.4118, 84.46875, 68.4174,
    60.60431, 61.6747, 58.62525, 57.46738, 58.04989, 59.21356, 61.04151,
    61.65593, 61.65002, 62.86916, 61.90791, 58.76103, 56.70959, 52.73343,
    48.83472, 46.98838, 47.58055, 48.39901, 47.84747, 45.61738, 42.88577,
    35.39835,
  78.06098, 81.72163, 84.7941, 85.1256, 86.96796, 92.84029, 89.44877,
    69.65573, 59.36187, 62.61201, 64.11179, 67.29469, 69.65215, 70.09549,
    69.36273, 67.7226, 62.73579, 57.03853, 53.69721, 49.44292, 45.81604,
    43.72315, 42.29848, 41.42032, 41.32667, 41.92644, 40.92753, 36.95753,
    33.02224, 28.96588,
  35.36404, 35.64212, 36.11514, 36.73563, 37.29877, 38.16624, 39.24092,
    40.49509, 42.03114, 44.07878, 47.11724, 48.51595, 46.49786, 48.17319,
    49.35834, 49.07475, 49.77304, 51.18373, 52.7709, 55.22277, 56.47779,
    55.00757, 55.652, 58.06718, 59.31432, 58.48817, 61.58102, 62.3348,
    47.04638, 42.08926,
  36.40867, 37.21778, 37.12213, 38.97055, 39.61444, 40.64569, 42.70509,
    44.88139, 47.38129, 50.27652, 53.77621, 57.7295, 60.4501, 59.69263,
    59.42078, 60.7007, 59.98798, 61.85191, 64.22684, 66.49635, 67.09562,
    66.57847, 66.64384, 69.41402, 72.36584, 67.07433, 58.91998, 62.05859,
    48.21394, 43.54241,
  37.51114, 39.07224, 40.80772, 42.78432, 44.70351, 46.747, 48.73488,
    50.91078, 53.39347, 55.83679, 58.30674, 61.33844, 64.14805, 66.98387,
    68.67365, 67.12272, 68.77438, 71.88364, 74.80838, 79.6875, 86.76926,
    92.42682, 91.77045, 87.58171, 83.88789, 78.48469, 70.83574, 60.18901,
    47.7356, 44.44102,
  44.60676, 47.31723, 50.61189, 54.00108, 56.89111, 59.58704, 60.59769,
    60.93493, 62.57472, 64.22724, 65.0322, 65.86804, 66.00772, 65.90619,
    70.14525, 72.55241, 70.18457, 69.01956, 74.43788, 80.69464, 89.56009,
    90.57985, 85.15837, 89.99525, 88.66242, 86.20261, 81.35537, 65.60902,
    51.13492, 43.2409,
  51.96186, 54.02859, 58.19488, 61.59929, 64.05682, 65.28362, 66.67967,
    68.15547, 71.03238, 73.14635, 73.36433, 75.55636, 77.13609, 77.73476,
    79.009, 79.97884, 76.85669, 72.00736, 74.12575, 80.60474, 81.32786,
    73.16171, 74.97397, 81.96132, 87.98328, 88.52997, 83.3166, 87.50069,
    77.99036, 52.0014,
  65.10148, 71.39003, 77.01958, 82.42873, 82.54517, 82.21961, 85.3362,
    86.32492, 86.98717, 89.27991, 93.81491, 103.1619, 111.8191, 107.8513,
    106.9633, 106.9506, 103.8254, 94.631, 83.03087, 80.98698, 73.23767,
    65.37698, 70.92937, 75.66626, 81.01849, 80.82769, 79.33047, 91.319,
    81.7648, 47.10749,
  75.90834, 81.4243, 86.33662, 91.01324, 92.01602, 93.90792, 100.4425,
    105.6909, 103.6203, 97.94135, 92.83008, 82.61209, 71.83635, 73.1272,
    75.12328, 78.16049, 79.23116, 75.50968, 69.85773, 70.92799, 68.36038,
    67.95765, 72.11216, 77.89197, 78.35429, 72.94424, 76.14743, 83.19147,
    69.79589, 40.62307,
  70.76659, 74.60432, 79.5702, 84.11292, 85.1991, 91.12384, 93.51479,
    77.76534, 70.38388, 71.79978, 69.82686, 67.83159, 67.25794, 69.77588,
    72.1375, 75.54689, 78.88052, 77.43864, 72.39407, 72.70744, 73.42287,
    76.20618, 81.14322, 83.38448, 79.13193, 77.34157, 83.76466, 80.715,
    59.60649, 42.34778,
  78.14102, 81.44877, 85.92841, 88.98589, 90.57974, 93.5955, 86.27829,
    87.58721, 93.0463, 96.29263, 97.56339, 97.34324, 99.62573, 108.2678,
    110.6998, 97.25014, 94.86463, 96.06673, 93.58161, 86.12818, 83.18436,
    89.84837, 96.77654, 93.62965, 83.41006, 87.11603, 84.5329, 69.61529,
    45.54138, 41.88748,
  106.3838, 113.6907, 108.4542, 110.4638, 111.3688, 104.5713, 88.74275,
    97.63556, 98.95023, 103.852, 109.3116, 114.7522, 110.3866, 105.4784,
    100.6062, 104.4792, 104.2097, 99.9652, 95.5712, 94.43076, 96.54613,
    91.73442, 85.42265, 76.96957, 80.62792, 88.05698, 77.24538, 52.55395,
    41.437, 39.32305,
  128.4064, 127.5435, 128.5169, 120.7304, 126.0585, 118.5688, 109.1306,
    111.2258, 111.321, 104.7154, 90.49318, 72.53067, 69.64409, 69.92899,
    70.57706, 72.806, 75.63631, 76.89322, 77.95433, 81.11327, 89.76833,
    84.2018, 70.16093, 67.05534, 71.04641, 67.24535, 51.92689, 42.28436,
    41.88874, 39.521,
  133.8823, 129.8295, 132.5814, 132.7197, 131.7882, 111.8106, 106.9547,
    97.70621, 87.57774, 77.50024, 72.51105, 69.59441, 72.74994, 73.61248,
    70.6656, 69.01212, 67.77782, 68.47308, 70.05093, 74.82877, 83.23952,
    80.27512, 69.3559, 77.13642, 77.88181, 60.52746, 44.10838, 47.12379,
    43.42415, 40.87247,
  140.8066, 140.6278, 142.1256, 142.1018, 140.0686, 134.986, 126.7692,
    117.6572, 122.9675, 103.5272, 97.93555, 92.24242, 98.84094, 100.7558,
    89.52048, 75.25798, 75.97845, 74.66402, 74.19312, 78.2281, 79.66487,
    72.36356, 65.93482, 61.56101, 60.05475, 53.19402, 45.01429, 46.3744,
    45.41223, 42.09952,
  129.7356, 129.9307, 129.8541, 129.078, 128.2711, 128.1858, 128.4238,
    128.2548, 125.8179, 125.6284, 126.1356, 124.9509, 126.012, 126.3919,
    114.8032, 93.82554, 88.83096, 92.31503, 93.92974, 85.10841, 72.72869,
    63.82828, 58.32374, 49.88112, 45.70586, 44.85442, 42.72929, 41.8649,
    42.24857, 41.33617,
  117.6276, 115.4841, 120.42, 124.2446, 126.7563, 127.7164, 129.1666,
    128.2975, 121.7535, 118.913, 110.8621, 103.4749, 104.1798, 106.056,
    103.0452, 99.14135, 89.49516, 85.58484, 85.25859, 78.01001, 61.11311,
    58.7717, 51.13075, 48.27243, 46.94921, 44.95488, 43.15057, 41.7168,
    40.60887, 40.00546,
  117.9968, 122.4296, 123.1973, 123.2992, 121.7063, 122.1068, 122.3707,
    112.1311, 98.91885, 92.63179, 90.40412, 84.3024, 79.95623, 86.82069,
    83.54165, 80.47357, 80.50748, 74.19144, 72.00909, 65.27522, 52.97663,
    54.09753, 49.46085, 47.80327, 46.99253, 45.33498, 43.07249, 42.00805,
    40.89704, 40.02758,
  99.83951, 97.87582, 99.12435, 101.1435, 102.4983, 103.7155, 103.5402,
    101.7483, 97.47153, 91.08571, 83.71975, 91.19697, 98.68054, 89.26492,
    82.14453, 76.54915, 71.48321, 68.38078, 69.73817, 65.06143, 52.54745,
    54.01648, 50.06499, 47.57054, 46.44862, 45.32007, 42.4334, 40.50191,
    40.24406, 39.87465,
  88.81033, 91.67551, 90.63919, 92.83575, 93.74152, 94.97002, 95.43523,
    95.72794, 96.2275, 96.2914, 104.8929, 111.5369, 106.699, 104.0729,
    96.39455, 86.43876, 76.76429, 75.103, 77.41518, 69.19321, 54.06742,
    52.74486, 49.50503, 47.79354, 44.75663, 43.10671, 42.00409, 39.85925,
    39.72503, 39.51783,
  99.63819, 92.06789, 80.54335, 74.21796, 74.59927, 74.17243, 75.81877,
    78.10338, 79.18963, 83.57593, 89.92681, 88.00558, 80.11478, 84.22097,
    86.48248, 89.16203, 96.03575, 101.1199, 97.54214, 84.16965, 64.49036,
    55.55875, 50.84248, 48.15055, 44.91603, 42.81012, 41.73031, 40.18143,
    39.6782, 39.52928,
  93.76769, 84.42633, 72.29039, 64.88995, 66.68695, 68.32451, 70.67281,
    72.73556, 75.75229, 80.92096, 80.11573, 68.80327, 68.5796, 68.61812,
    68.37148, 69.13123, 74.36638, 81.44818, 84.18779, 81.64583, 73.21187,
    63.46661, 54.93139, 50.98368, 47.49847, 43.78222, 41.91616, 40.42023,
    39.62928, 39.52808,
  86.83037, 77.39815, 67.27255, 61.57224, 62.97282, 63.9644, 64.57131,
    64.72924, 65.74981, 67.4278, 62.02897, 55.24325, 59.74588, 59.82441,
    58.53408, 57.97173, 60.06651, 63.08688, 66.65085, 67.76356, 67.97124,
    68.01114, 62.12948, 55.47783, 49.92429, 45.06023, 41.85207, 40.39499,
    39.64132, 39.54789,
  85.31872, 77.08684, 68.21268, 64.0065, 63.76923, 60.69094, 60.54195,
    59.50788, 61.65585, 61.02112, 53.34968, 49.63059, 52.90133, 53.43884,
    53.03196, 53.65239, 54.41195, 55.84238, 58.80688, 60.62407, 61.34352,
    61.67904, 62.1512, 61.37464, 55.21621, 46.65999, 42.50117, 41.25998,
    39.92038, 39.50471,
  86.89708, 82.72876, 72.19096, 68.62431, 70.71139, 69.799, 66.58096,
    61.3672, 60.67148, 57.57363, 51.14268, 53.11617, 55.11067, 56.35343,
    55.83698, 57.41032, 58.01718, 55.81448, 56.04582, 57.06292, 57.34491,
    57.22072, 56.88906, 59.07991, 59.82475, 52.32786, 45.45929, 43.82114,
    41.6221, 39.72437,
  95.68742, 91.86843, 87.8575, 84.6088, 84.5997, 82.19488, 81.9429, 79.94954,
    79.16791, 71.51447, 64.10673, 68.57184, 70.91901, 72.11681, 70.46368,
    69.65749, 68.57785, 65.01619, 61.32442, 60.21187, 59.00712, 57.85524,
    56.98052, 56.93349, 58.9128, 59.29175, 53.45378, 46.65971, 44.26583,
    40.9668,
  94.39962, 91.13418, 81.12471, 78.89503, 78.76398, 77.54788, 77.9006,
    80.2187, 84.22354, 75.78482, 67.73213, 72.19318, 74.42613, 75.48741,
    74.65096, 73.60493, 70.56006, 68.19926, 65.8374, 62.50048, 60.86373,
    59.14706, 56.28092, 54.67005, 55.78238, 58.82726, 59.15646, 52.04037,
    47.29156, 43.22924,
  101.6872, 98.49207, 92.53717, 85.21619, 81.11845, 79.79005, 83.6776,
    86.90592, 82.69974, 74.51839, 73.51702, 75.63529, 77.32231, 75.59925,
    73.58085, 73.15756, 71.83172, 70.62941, 70.28161, 68.10784, 66.47639,
    64.46521, 60.28002, 57.46086, 57.85726, 59.43052, 60.82246, 54.11486,
    44.99134, 41.88841,
  102.1002, 96.71642, 88.21678, 83.63188, 79.97987, 75.8145, 80.25209,
    80.29004, 74.81763, 72.5158, 76.12496, 78.71925, 79.38269, 77.76805,
    76.42496, 75.1073, 73.65167, 73.15102, 73.53762, 73.24001, 73.16305,
    73.74696, 71.80494, 67.87008, 67.01814, 68.40506, 70.38182, 63.17208,
    47.66461, 40.24035,
  101.7242, 95.69102, 91.88388, 90.62798, 89.22769, 85.2995, 83.02573,
    77.57645, 70.53085, 72.40772, 73.85301, 75.83822, 77.1208, 76.81467,
    76.38185, 74.81944, 71.89819, 71.00778, 72.67125, 73.77404, 71.25182,
    66.85191, 62.72324, 61.12815, 62.11975, 63.7779, 65.15966, 66.58298,
    59.22698, 44.18422,
  86.93336, 84.38041, 87.86765, 91.32818, 94.17617, 96.17216, 86.06936,
    71.9119, 66.53882, 66.60927, 64.32924, 63.91287, 64.51311, 64.93188,
    65.6115, 65.18115, 63.40897, 61.99229, 59.77821, 56.86067, 55.6074,
    54.05436, 51.41853, 49.9001, 51.08327, 52.37222, 52.37135, 50.70975,
    50.3066, 45.54316,
  76.81414, 78.31553, 77.16844, 75.75163, 79.59332, 86.27385, 84.78278,
    69.24216, 62.16123, 64.88265, 66.14053, 67.66948, 67.51819, 65.17212,
    62.05746, 58.68097, 53.40778, 49.18678, 48.51604, 47.4815, 45.70942,
    45.96542, 46.0712, 46.0862, 46.64667, 47.84399, 47.78149, 45.08302,
    42.07325, 39.54017,
  47.82195, 48.96451, 49.74622, 50.66551, 51.17991, 51.79863, 52.51805,
    53.17011, 53.83113, 54.61251, 55.79035, 55.69858, 53.06302, 52.99496,
    52.6299, 50.9961, 50.19394, 50.10336, 50.19333, 50.87413, 50.75797,
    48.95419, 49.25631, 51.216, 52.43698, 51.35733, 52.85871, 54.09566,
    43.62701, 39.87868,
  55.01907, 56.39921, 56.33676, 57.84034, 58.08486, 58.43612, 59.44259,
    60.28434, 61.11417, 62.01768, 63.28501, 64.76864, 65.28094, 63.43257,
    61.90982, 61.36343, 59.80545, 60.05402, 60.83127, 61.46685, 60.82207,
    59.73619, 59.33574, 61.66792, 64.06135, 58.30354, 50.65537, 53.54974,
    44.46824, 40.86484,
  57.66639, 58.83102, 59.44258, 60.18754, 60.64486, 61.15384, 61.62971,
    62.10226, 62.66486, 63.23322, 63.91753, 65.14215, 66.2562, 67.43549,
    67.84598, 65.75204, 65.90953, 67.46291, 69.24341, 72.29129, 77.33952,
    81.71031, 80.86002, 76.55936, 73.14835, 68.21577, 60.72021, 52.39789,
    43.92075, 41.54581,
  63.63942, 64.92834, 66.0986, 67.35457, 68.1726, 68.93029, 68.60027,
    67.67017, 67.56378, 67.41836, 66.98031, 67.14567, 66.72484, 65.86009,
    67.78859, 68.33202, 65.57126, 64.2697, 67.71577, 71.82677, 78.0146,
    77.83965, 72.24182, 75.4161, 74.06151, 72.14923, 70.01625, 57.64054,
    46.43615, 40.70896,
  70.8512, 71.09959, 72.41294, 73.32393, 73.60709, 73.45531, 73.62302,
    73.47784, 74.28149, 74.77088, 74.58778, 76.12891, 76.72748, 75.66288,
    75.59093, 75.58838, 72.06899, 67.42914, 67.77848, 71.88546, 71.21805,
    63.03632, 63.72121, 68.65754, 73.1577, 74.30517, 71.72549, 75.71698,
    68.0087, 48.08431,
  75.02136, 78.03049, 80.55058, 82.82297, 81.75004, 81.33344, 83.73311,
    84.00299, 82.95174, 83.22885, 85.92725, 93.38874, 100.1899, 96.42404,
    95.96434, 96.01469, 92.27592, 84.59653, 74.90506, 71.81165, 64.46464,
    56.5038, 60.75978, 64.20233, 68.23833, 68.89095, 68.63181, 78.77283,
    73.14942, 43.72147,
  77.57655, 81.65314, 84.93154, 87.94232, 88.56885, 90.94639, 96.96692,
    101.0535, 98.88213, 93.05161, 88.43943, 79.9796, 69.79585, 69.6637,
    70.27209, 71.86238, 71.90199, 68.20854, 63.81005, 63.4118, 60.20478,
    58.59207, 61.22377, 65.01699, 65.43899, 62.46581, 65.97157, 71.6401,
    60.64587, 38.46384,
  82.99533, 86.76029, 89.9792, 92.98892, 93.93255, 99.05258, 101.2486,
    86.81403, 79.18851, 78.74347, 75.38997, 72.01156, 69.38101, 68.79994,
    68.31512, 69.18392, 71.02747, 69.65849, 65.18896, 63.91908, 63.13094,
    64.5565, 67.8453, 69.46671, 66.75301, 66.29551, 71.88051, 69.57629,
    52.5458, 39.49129,
  91.6555, 92.79102, 93.28677, 93.68942, 93.97778, 94.68466, 86.17188,
    85.12059, 87.46107, 87.58684, 86.81932, 85.41382, 85.06721, 89.28411,
    90.4709, 82.26408, 81.04395, 81.83511, 78.93015, 72.33138, 68.75428,
    72.36648, 77.56365, 76.12324, 70.13359, 73.77819, 73.21764, 61.46944,
    41.75716, 39.42253,
  105.3259, 107.1051, 99.61959, 98.63621, 97.69597, 90.68443, 75.71352,
    80.78925, 79.74803, 81.36739, 83.16362, 86.18109, 84.09186, 82.27188,
    79.86882, 83.00674, 83.75513, 81.71922, 78.08644, 76.51434, 76.69056,
    72.82265, 69.05687, 64.27689, 68.18559, 75.84523, 68.11339, 47.63432,
    39.26414, 37.8636,
  127.4363, 126.8148, 124.5533, 109.7867, 109.9567, 98.76632, 90.088,
    89.74747, 89.22862, 85.91081, 75.50286, 62.94918, 61.24345, 61.44557,
    62.1633, 63.35626, 64.70909, 65.25252, 65.7907, 67.73553, 73.25542,
    69.78827, 61.05056, 59.90611, 63.85284, 61.44308, 48.20542, 39.86576,
    39.72618, 37.97643,
  135.38, 132.261, 133.5831, 132.5959, 129.506, 110.7765, 102.7521, 92.78275,
    84.92895, 78.23161, 73.30341, 69.08162, 70.45766, 69.7924, 65.01308,
    63.0733, 61.26277, 60.59227, 60.55711, 63.21869, 68.60523, 67.11353,
    60.75144, 67.45367, 69.82693, 56.41014, 41.4007, 43.97754, 40.79778,
    38.94314,
  134.7743, 135.7905, 136.9042, 136.5435, 134.9692, 131.6276, 125.0101,
    112.3711, 114.708, 100.0114, 94.53506, 88.19807, 91.17042, 92.25136,
    82.05621, 67.82436, 67.79205, 65.88692, 63.86839, 64.96599, 65.71794,
    61.44055, 57.51868, 54.63042, 54.12427, 49.37057, 42.42067, 43.30983,
    42.42381, 39.93204,
  114.7652, 115.6094, 112.0555, 110.9662, 109.618, 117.2305, 125.2713,
    124.2902, 109.836, 111.7062, 115.0027, 110.5429, 109.1388, 107.1108,
    97.32616, 82.80861, 75.54359, 78.35123, 78.73399, 71.29663, 62.70128,
    56.20144, 51.63127, 45.48523, 42.35709, 42.16692, 40.66197, 39.87916,
    40.05751, 39.29219,
  87.30331, 84.29982, 86.36417, 87.33858, 89.13232, 91.10648, 95.57374,
    95.52171, 90.13595, 89.36081, 87.23445, 82.35884, 83.79067, 87.60678,
    86.94228, 83.65082, 76.91592, 72.52362, 70.70537, 65.50179, 53.68547,
    51.83376, 46.08614, 43.65023, 43.07518, 42.01483, 40.82014, 39.65376,
    38.85611, 38.37055,
  86.60514, 89.41719, 90.12739, 89.71759, 88.98059, 90.95594, 93.15207,
    87.5943, 81.80721, 77.33143, 75.32187, 72.34254, 70.00356, 74.12446,
    71.40332, 69.80949, 69.70222, 64.13431, 60.779, 55.73357, 48.5122,
    48.48943, 44.69017, 43.44036, 43.00634, 42.18367, 40.81468, 39.87017,
    38.98784, 38.34932,
  77.63158, 77.01036, 78.10548, 80.3131, 82.44355, 84.19315, 86.09419,
    88.08629, 85.67484, 81.16815, 76.27137, 80.97546, 85.32786, 79.29644,
    72.19487, 67.84311, 63.76511, 60.78252, 59.61315, 55.96416, 47.86496,
    48.33213, 45.13185, 43.39116, 42.77413, 42.16604, 40.33316, 38.81732,
    38.54369, 38.25368,
  72.36187, 73.25692, 72.28104, 74.55495, 76.69928, 79.07879, 80.99913,
    83.33878, 84.97906, 84.36026, 88.95981, 92.93396, 90.83968, 88.84723,
    82.88539, 76.72606, 71.27277, 68.70599, 67.57361, 60.0066, 49.30668,
    47.2166, 44.93577, 43.68619, 41.85625, 40.82421, 39.95552, 38.33167,
    38.13561, 37.96061,
  79.12965, 73.87781, 65.96323, 62.99266, 65.50893, 66.48737, 68.35376,
    70.13225, 70.56384, 72.77746, 76.82816, 75.45936, 70.10371, 72.3055,
    72.74279, 74.72669, 80.19589, 83.99415, 81.13635, 71.57715, 57.71178,
    49.87291, 46.04048, 44.20169, 42.08389, 40.56675, 39.6601, 38.46599,
    38.09789, 37.97367,
  72.97997, 68.35455, 60.70013, 56.26849, 58.13214, 59.25784, 60.74586,
    62.20955, 64.41441, 68.58488, 68.78578, 62.61722, 62.42908, 61.04059,
    59.67339, 59.54461, 62.82889, 67.80757, 69.34447, 67.907, 62.26266,
    54.86139, 49.04332, 46.24354, 43.86851, 41.25239, 39.85094, 38.66833,
    38.07156, 37.97882,
  70.95148, 66.93153, 58.88375, 54.75071, 55.43909, 56.15163, 57.28362,
    58.56638, 60.60097, 62.55534, 59.73011, 56.0192, 58.64398, 57.903,
    55.92157, 54.6784, 55.18489, 56.44395, 58.1382, 58.10962, 57.64074,
    57.52782, 53.68144, 49.38924, 45.53547, 42.05788, 39.94143, 38.72469,
    38.07435, 37.99013,
  75.01424, 71.94907, 64.91373, 61.53811, 61.53837, 59.99091, 60.24538,
    60.20559, 62.29226, 62.10117, 57.15736, 54.62623, 55.85957, 55.38624,
    54.161, 53.61471, 52.82515, 52.58978, 53.48606, 53.79648, 53.58461,
    53.24847, 53.28667, 52.51223, 48.46227, 43.03388, 40.53574, 39.40042,
    38.26445, 37.94069,
  82.23284, 81.94337, 74.19605, 71.57453, 73.84546, 73.8903, 71.64846,
    67.97777, 67.48434, 65.16409, 60.34934, 60.61844, 60.60994, 60.0397,
    58.11926, 57.48136, 56.15595, 53.28831, 52.20938, 51.70951, 50.98987,
    50.42511, 49.88286, 51.12728, 51.61253, 46.99247, 42.69839, 41.26009,
    39.52138, 38.11889,
  87.97632, 87.48207, 82.10944, 80.29639, 80.61008, 79.86668, 80.13824,
    78.94576, 79.8914, 74.85095, 69.91861, 71.68599, 72.26457, 71.92996,
    69.38622, 66.89609, 64.49174, 60.53391, 56.31622, 54.11674, 52.34491,
    51.09593, 50.20718, 49.90982, 51.43903, 52.04801, 48.19663, 43.34818,
    41.52587, 39.10813,
  90.25603, 86.24471, 78.96331, 76.29959, 76.02143, 75.32342, 76.50953,
    79.70829, 83.407, 77.82333, 71.43785, 72.89407, 73.37534, 73.54889,
    71.73551, 69.71088, 67.0327, 64.2562, 60.59336, 56.9901, 55.11439,
    53.2859, 50.66119, 49.3596, 50.42785, 52.52918, 52.25476, 47.08404,
    43.70356, 40.72948,
  94.28912, 91.5871, 85.94734, 80.13958, 76.96852, 75.72835, 79.48281,
    83.63609, 82.40736, 76.58335, 74.77142, 74.46719, 74.74449, 73.3513,
    70.65747, 69.07016, 67.85422, 66.14867, 63.78871, 60.93723, 59.7566,
    58.16694, 54.33833, 51.86915, 52.02159, 52.38015, 52.5225, 48.18929,
    42.0978, 39.78284,
  92.94958, 89.12743, 82.65862, 78.37309, 75.068, 72.26137, 75.66502,
    76.6339, 73.7721, 71.67722, 72.78542, 73.13202, 72.93065, 71.97354,
    70.18433, 68.72325, 67.56033, 66.61955, 65.08826, 63.57214, 63.74787,
    64.27446, 62.02019, 59.0294, 58.10386, 57.9039, 57.84178, 53.60559,
    43.72439, 38.66464,
  85.55856, 83.42355, 79.79615, 78.42401, 77.45474, 74.12207, 71.55031,
    67.82716, 63.40404, 63.91022, 64.6969, 65.93632, 67.14134, 67.41499,
    66.94509, 65.56699, 63.77563, 62.99294, 62.98908, 62.68742, 61.20164,
    58.65808, 55.90778, 54.78674, 55.27898, 55.63957, 55.44907, 55.86326,
    51.07266, 41.38089,
  68.31994, 68.1295, 69.3968, 70.29384, 72.52254, 74.23325, 68.7581,
    59.07502, 55.91827, 56.84544, 56.3441, 56.70774, 57.59211, 58.20832,
    58.4241, 57.75435, 56.05936, 54.79223, 52.89376, 50.78732, 50.20242,
    49.50133, 47.89356, 47.05791, 47.96452, 48.69169, 47.90951, 46.13202,
    45.50638, 42.11415,
  55.19194, 55.85413, 55.35078, 54.80009, 57.38092, 62.46367, 62.87793,
    53.90964, 49.7501, 52.12204, 53.69101, 55.18225, 55.65958, 54.51284,
    52.81847, 51.07788, 47.59471, 44.87449, 44.53361, 43.78642, 42.78782,
    43.17897, 43.46917, 43.4997, 43.84668, 44.66946, 44.31035, 42.03869,
    39.85387, 38.03271,
  43.55996, 43.71905, 43.82224, 43.98236, 44.08247, 44.25416, 44.48941,
    44.80857, 45.17625, 45.797, 46.8146, 46.70246, 44.81107, 45.33858,
    45.70957, 45.41821, 45.66378, 46.23266, 46.83118, 47.88382, 48.40603,
    47.454, 48.15388, 50.2328, 51.75507, 51.14773, 52.17873, 52.99985,
    44.79484, 42.15236,
  48.60357, 48.77774, 48.16305, 48.59289, 48.23445, 48.02552, 48.34029,
    48.54773, 48.84217, 49.29855, 50.03156, 50.87051, 51.25325, 50.24678,
    49.73257, 50.36702, 49.96181, 50.85555, 51.86662, 52.67097, 52.77285,
    52.84478, 54.07323, 57.70224, 60.75645, 56.14744, 49.40641, 52.40733,
    45.37588, 42.82424,
  51.61368, 51.7365, 51.72165, 51.79572, 51.86007, 52.11262, 52.4107,
    52.81135, 53.24957, 53.72607, 54.35093, 55.25141, 56.27909, 57.54265,
    58.32608, 57.44907, 58.38317, 60.19035, 61.74719, 64.32933, 68.88059,
    73.62667, 74.14986, 71.07721, 68.47084, 64.06966, 58.10507, 51.90565,
    45.31758, 43.5327,
  55.48279, 55.95881, 56.55794, 57.29536, 57.7935, 58.42533, 58.40348,
    58.24211, 58.64322, 59.07454, 59.1889, 59.55203, 59.49126, 59.076,
    61.0218, 62.18863, 61.08493, 60.86162, 63.97639, 67.74297, 73.09383,
    73.12847, 67.71809, 70.04817, 67.7472, 66.04366, 64.49535, 54.73312,
    46.14331, 42.55197,
  58.66778, 58.16175, 58.9319, 59.48931, 59.68785, 59.52815, 59.77896,
    60.03814, 61.0568, 61.67812, 61.54581, 62.86655, 63.63897, 63.66321,
    64.46664, 65.88404, 65.17725, 63.42237, 65.64859, 70.27626, 70.0057,
    62.03058, 61.67308, 65.98605, 69.05209, 69.03976, 67.09964, 71.53268,
    67.04351, 49.74847,
  65.05363, 67.12311, 69.10147, 71.14492, 70.79993, 70.83676, 73.11464,
    74.15365, 74.92656, 76.64229, 80.29294, 88.24445, 95.14554, 91.60815,
    92.06131, 93.46143, 90.58958, 83.51904, 75.56178, 72.67251, 65.48168,
    58.11202, 62.1747, 65.42828, 69.15264, 69.70753, 70.21722, 79.53807,
    73.39782, 46.4933,
  70.83356, 73.63152, 76.20718, 78.78748, 79.83595, 82.66039, 89.05865,
    94.20264, 93.4626, 88.57689, 84.60794, 77.07252, 68.18343, 69.0414,
    70.42151, 71.92566, 72.25119, 68.72399, 64.06396, 62.95987, 59.3405,
    57.80331, 60.65308, 64.31308, 65.29005, 63.06316, 66.70609, 72.20044,
    61.33863, 40.99158,
  69.32883, 71.41893, 73.61015, 75.84406, 76.77023, 81.44114, 83.70828,
    70.99135, 63.82793, 63.72751, 61.23019, 58.5987, 57.20064, 58.25869,
    59.72583, 62.23412, 64.67257, 64.07645, 61.00973, 60.45062, 59.84282,
    60.93765, 64.06934, 66.68156, 65.9912, 66.80146, 72.65579, 70.06086,
    54.13654, 41.36773,
  74.56355, 75.69717, 76.74651, 77.49458, 78.96097, 80.02951, 71.71997,
    69.87794, 71.83919, 72.17062, 72.19846, 71.87421, 72.78328, 77.30205,
    79.66922, 74.37714, 75.2214, 77.2386, 75.57497, 70.23892, 67.22073,
    70.03687, 74.20889, 73.51687, 69.73088, 74.1776, 74.24377, 62.88256,
    43.73532, 41.93793,
  85.86649, 89.52397, 85.0285, 86.21423, 88.07384, 82.7485, 68.51413,
    73.92558, 73.90696, 76.45163, 79.08975, 82.77028, 81.25407, 79.72618,
    77.86096, 80.03122, 80.50803, 79.29008, 76.89626, 75.72546, 75.50806,
    72.20894, 69.27982, 65.70878, 69.81109, 76.63422, 68.9157, 49.73501,
    41.64059, 40.73329,
  108.6189, 106.9403, 102.9337, 92.58015, 94.65263, 85.46547, 76.49679,
    78.6831, 79.81111, 77.53467, 70.0225, 60.73679, 59.61737, 60.33241,
    61.09038, 62.23286, 63.50896, 63.87676, 64.21449, 65.86635, 70.2664,
    67.26387, 60.11597, 59.17233, 63.90236, 62.80096, 50.31339, 41.80508,
    42.24619, 40.75587,
  117.1868, 113.0652, 116.2119, 115.5975, 105.0293, 84.71506, 81.61372,
    74.1431, 68.08665, 65.49859, 62.0915, 60.12201, 62.07546, 61.92679,
    59.73163, 59.73191, 58.98099, 59.29671, 59.49988, 61.67832, 66.40278,
    65.78499, 60.30724, 66.39796, 68.85442, 56.6808, 42.64228, 45.02392,
    42.65707, 41.46708,
  123.5032, 123.9943, 124.546, 123.1417, 120.0481, 115.1699, 101.3106,
    86.57867, 91.26717, 80.65971, 76.14896, 72.67644, 76.38137, 78.21893,
    72.05612, 62.03894, 62.70805, 62.37243, 61.95543, 63.70042, 65.65462,
    63.61971, 60.60462, 57.74149, 56.12949, 50.7627, 44.18785, 45.05132,
    44.10888, 42.34713,
  114.7004, 114.9879, 114.1225, 111.6961, 109.1327, 110.1994, 110.3555,
    108.7753, 99.35655, 98.74724, 102.2166, 97.93537, 95.97687, 96.02997,
    89.51745, 75.71239, 71.80008, 74.78194, 75.87239, 69.73962, 63.01954,
    58.21864, 53.84365, 47.77814, 44.7574, 44.26323, 42.97821, 42.47136,
    42.54581, 41.88981,
  86.27029, 82.9693, 84.58641, 84.57774, 85.86821, 89.12221, 94.66893,
    93.00601, 87.48415, 86.45857, 82.80403, 78.60075, 80.39137, 83.29868,
    83.04001, 81.7578, 74.50623, 70.57639, 68.48878, 64.32726, 55.43293,
    52.853, 47.1962, 44.81541, 44.56075, 43.88177, 42.82236, 41.98856,
    41.5043, 41.13453,
  76.78059, 78.87583, 79.54388, 78.83406, 77.50312, 78.37704, 80.49542,
    77.7411, 72.70284, 69.31566, 68.62398, 66.53296, 65.32995, 69.04665,
    67.41902, 66.52271, 66.64172, 62.17158, 59.40638, 55.35084, 48.93246,
    49.00114, 45.64487, 44.52988, 44.40907, 44.00876, 42.91026, 42.16271,
    41.51348, 41.09731,
  67.45598, 66.1583, 66.29138, 67.12419, 67.98053, 68.69485, 69.90868,
    71.44427, 70.15437, 67.66943, 64.14898, 68.166, 72.43159, 68.95103,
    64.6888, 62.35668, 59.78271, 58.08307, 58.05699, 55.46159, 49.14806,
    49.22712, 46.25069, 44.74979, 44.41148, 44.11852, 42.62714, 41.46543,
    41.20111, 40.98964,
  64.45577, 64.96591, 63.83484, 64.88909, 65.79523, 67.11172, 68.3261,
    69.85287, 70.96477, 70.35818, 74.06353, 77.28695, 76.01761, 74.84691,
    69.84747, 65.49739, 61.22234, 60.34805, 60.92511, 56.44215, 49.25611,
    48.15549, 46.2905, 45.27419, 43.89982, 43.06926, 42.31189, 41.04294,
    40.91132, 40.80686,
  73.53152, 69.00754, 62.25193, 59.26128, 60.98043, 61.42969, 62.54033,
    63.8399, 64.185, 66.2206, 69.93709, 69.47611, 64.90093, 66.33765,
    66.2334, 67.85507, 72.22415, 75.49463, 73.27371, 65.88535, 55.69431,
    49.70452, 46.80156, 45.66143, 43.97712, 42.7625, 42.05045, 41.17875,
    40.88028, 40.78793,
  70.17031, 65.98701, 59.78579, 55.96503, 57.42651, 58.13867, 59.12824,
    60.14993, 61.96875, 65.2987, 66.019, 61.85543, 61.79669, 60.78662,
    59.56767, 59.62114, 62.14681, 65.60304, 65.5125, 63.15541, 58.45895,
    52.61321, 48.24256, 46.96429, 45.27592, 43.2769, 42.23195, 41.3017,
    40.8486, 40.80288,
  66.11996, 62.53387, 56.04268, 52.57617, 53.20357, 53.65246, 54.40139,
    55.36677, 57.10506, 58.84003, 56.96884, 54.2464, 56.53712, 56.31874,
    54.97703, 54.33405, 55.05822, 56.01566, 56.60196, 55.83067, 55.09027,
    54.60538, 51.70665, 48.8523, 46.3254, 43.93716, 42.27146, 41.30415,
    40.84774, 40.82085,
  64.54343, 61.54596, 55.25589, 52.4307, 52.76562, 51.90617, 52.66219,
    53.28064, 55.41203, 55.76166, 52.24576, 50.43742, 52.03353, 52.33206,
    51.95902, 52.29126, 52.65457, 53.19352, 53.81779, 54.01628, 53.8925,
    53.38043, 53.04207, 51.51896, 48.19221, 44.58445, 42.6895, 41.75423,
    40.96323, 40.79802,
  66.89664, 65.72919, 58.64912, 56.04979, 57.7633, 57.8027, 56.89712,
    55.01819, 55.11892, 53.7955, 50.46683, 51.06931, 51.99348, 52.73885,
    52.424, 53.04172, 53.4654, 52.50303, 51.97182, 51.75129, 51.45792,
    51.04744, 50.3171, 50.28589, 50.229, 47.06269, 44.12578, 43.11082,
    41.82642, 40.90549,
  73.31458, 72.94545, 67.91396, 65.65034, 65.64169, 64.43129, 64.70168,
    64.16829, 65.32019, 62.40841, 59.09083, 60.6902, 61.86578, 62.59949,
    61.50751, 60.62475, 60.11252, 57.77515, 54.60102, 53.03622, 51.86585,
    51.25389, 50.48575, 49.71515, 50.60255, 51.06086, 48.29125, 44.59261,
    43.13472, 41.54538,
  76.08363, 72.6051, 66.11787, 63.39405, 63.41703, 62.96433, 64.01495,
    66.5938, 69.68405, 66.2429, 62.30071, 64.26283, 65.6021, 66.05621,
    65.17503, 64.94672, 63.60749, 61.59125, 58.79256, 56.33302, 54.67856,
    53.13658, 51.10275, 50.00947, 50.98113, 52.36727, 51.69339, 47.82496,
    45.27373, 42.90673,
  79.07709, 76.98676, 70.95693, 65.76437, 64.44253, 64.06163, 66.98588,
    70.2578, 69.55481, 65.55147, 64.5984, 65.70918, 66.97787, 65.83128,
    64.04604, 64.16435, 63.69377, 62.312, 60.67125, 58.65643, 57.09287,
    55.14862, 52.32267, 51.00945, 51.55434, 51.53967, 51.49859, 48.68745,
    44.25929, 42.25893,
  79.52465, 76.74546, 71.14865, 67.37271, 65.73286, 64.11768, 67.10614,
    68.29953, 66.6814, 64.85516, 65.92766, 67.19324, 67.8941, 66.87016,
    65.50461, 65.16676, 64.68889, 63.82729, 62.6836, 61.81463, 61.38628,
    61.17869, 59.47725, 57.52806, 56.92788, 56.09617, 55.60779, 52.51834,
    45.15141, 41.27853,
  77.41258, 75.60565, 72.87228, 71.97369, 72.21382, 70.39497, 69.4167,
    67.36565, 64.03148, 64.36849, 65.24259, 66.99292, 68.4621, 68.39644,
    67.83405, 66.72495, 65.52129, 64.99929, 64.99339, 64.68409, 62.82674,
    59.88421, 57.28395, 56.41409, 56.41357, 56.01886, 55.24674, 55.08077,
    50.90971, 43.16114,
  65.81715, 66.15778, 67.15256, 68.05811, 70.09881, 71.37867, 67.56256,
    60.78165, 58.22152, 58.3955, 57.78321, 58.36744, 59.77822, 61.07137,
    61.77992, 61.18929, 59.54349, 58.15831, 56.17738, 54.22065, 53.1513,
    51.96151, 50.3935, 49.60291, 50.15147, 50.51414, 49.71602, 47.8106,
    46.79234, 44.04489,
  59.57113, 60.30088, 60.50843, 60.30558, 62.63852, 66.85335, 66.97309,
    59.67007, 56.33631, 57.79301, 58.50533, 59.64569, 59.92607, 59.07682,
    57.82296, 55.82316, 52.34241, 49.6059, 48.89639, 47.8264, 46.81394,
    46.86985, 47.00618, 46.93284, 47.03284, 47.51192, 46.79876, 44.43449,
    42.56336, 40.94181,
  43.87958, 43.88844, 43.95703, 44.00638, 44.01741, 44.15223, 44.38271,
    44.6808, 45.00959, 45.45716, 46.27246, 46.19001, 44.67837, 44.9617,
    45.07827, 44.64197, 44.68975, 44.98484, 45.39674, 46.21387, 46.59209,
    45.94848, 46.50461, 48.37629, 50.18751, 50.48885, 51.9782, 53.26093,
    47.08939, 44.84825,
  45.05373, 45.15627, 44.80798, 45.22449, 44.99876, 44.98515, 45.36993,
    45.74476, 46.17763, 46.61303, 47.11357, 47.57717, 47.61995, 46.71677,
    46.20168, 46.55128, 46.09224, 46.75689, 47.80557, 48.78374, 49.02502,
    49.55097, 51.71947, 56.50978, 60.5883, 56.53936, 50.95874, 53.79591,
    47.91054, 45.56883,
  44.77697, 44.74548, 44.79976, 44.84826, 44.87167, 45.10498, 45.39468,
    45.72401, 46.10885, 46.49374, 46.9473, 47.59815, 48.32819, 49.233,
    49.95006, 49.69304, 50.80054, 52.89463, 54.95657, 58.09926, 63.05779,
    68.98111, 71.36713, 69.95017, 68.15075, 63.22406, 58.39785, 53.3014,
    47.95079, 46.19442,
  46.1967, 46.69843, 47.5247, 48.42013, 49.03762, 49.80241, 50.10307,
    50.13023, 50.64689, 51.26723, 51.791, 52.72009, 53.39217, 53.78333,
    56.2239, 58.3056, 58.74507, 59.76963, 63.74244, 68.48564, 74.48818,
    74.55891, 68.83739, 69.50932, 66.68597, 65.20415, 63.72857, 55.3745,
    47.71064, 45.07954,
  49.91174, 49.89434, 50.92354, 51.71258, 51.99784, 51.90251, 51.88816,
    51.83262, 52.43145, 52.75927, 52.65399, 53.84475, 55.30314, 56.94189,
    59.09, 61.73796, 62.67759, 62.85842, 66.2826, 71.08434, 70.83969,
    63.13266, 61.22313, 65.03391, 67.32909, 67.00377, 65.79839, 70.73344,
    67.34879, 52.04321,
  51.07097, 52.01592, 53.46174, 54.8359, 54.29017, 54.03838, 55.87053,
    57.49383, 59.79471, 63.37583, 68.6521, 78.47301, 87.47578, 86.00478,
    88.23163, 90.06838, 88.20026, 83.77929, 77.55042, 74.4244, 67.01336,
    59.73421, 64.10018, 67.81877, 71.9203, 72.58646, 73.06082, 82.48107,
    76.63026, 49.66409,
  56.11189, 59.10965, 62.33786, 65.8126, 68.59268, 74.06485, 83.91508,
    92.80646, 93.82671, 93.63956, 93.73619, 88.86313, 81.39621, 81.02936,
    80.99243, 81.01491, 80.52115, 75.90308, 70.27911, 68.40797, 64.47346,
    63.05963, 66.18907, 69.63033, 70.88343, 68.88385, 71.6214, 76.27238,
    64.16544, 43.81046,
  67.08877, 72.11913, 76.5682, 81.11186, 84.43927, 91.81618, 94.53791,
    85.72752, 77.19006, 75.1393, 70.87073, 66.41133, 63.47263, 63.2981,
    63.69028, 65.24702, 66.44892, 65.37378, 63.11002, 62.9359, 62.52126,
    63.56469, 66.42435, 68.61422, 67.89761, 68.67926, 73.92202, 71.4464,
    56.4597, 43.79585,
  74.16699, 77.03906, 78.59363, 79.24959, 80.79868, 80.81684, 70.8628,
    65.39355, 64.95097, 63.95469, 63.07884, 63.09972, 64.70023, 69.13632,
    71.6273, 67.80865, 68.91272, 71.32402, 71.06757, 68.08473, 66.61538,
    70.21539, 74.43915, 73.95264, 71.72133, 76.67342, 77.30798, 65.38647,
    46.4787, 44.54479,
  78.92377, 82.30079, 78.05956, 77.97724, 78.89091, 73.7766, 59.76129,
    64.67883, 66.03122, 69.70906, 73.86739, 78.06143, 78.13492, 77.33332,
    75.7316, 77.45483, 78.75186, 78.44114, 77.03137, 76.70246, 76.88953,
    74.62743, 72.14912, 68.66917, 72.83468, 80.03231, 72.99895, 52.97874,
    44.10695, 43.77514,
  79.46662, 80.23843, 81.06544, 80.82565, 84.67828, 78.81703, 72.16045,
    76.93709, 81.09779, 82.25987, 76.17894, 67.31861, 65.83396, 66.14472,
    66.62025, 67.86615, 68.99465, 69.08622, 69.33154, 71.30009, 74.73729,
    71.23077, 64.47158, 63.48627, 69.2411, 68.73682, 54.71844, 44.40991,
    44.88935, 43.66092,
  87.46776, 82.47421, 90.30317, 95.37804, 90.27561, 79.449, 81.23452,
    75.12874, 69.66267, 68.37398, 64.23502, 61.58054, 63.85121, 64.21148,
    62.43345, 62.97885, 62.43819, 62.68463, 63.04755, 65.11755, 69.25848,
    68.53922, 64.00605, 69.59968, 71.98335, 59.78273, 45.03262, 47.10742,
    45.27226, 44.2044,
  102.81, 105.2824, 107.6005, 107.3836, 105.398, 101.9527, 88.3353, 75.9257,
    81.07742, 73.13287, 69.74458, 68.83528, 73.42769, 75.51755, 70.25744,
    61.45123, 62.9059, 63.21907, 63.82321, 66.35067, 69.6039, 69.29017,
    66.65134, 63.28868, 60.28468, 53.75859, 46.51394, 47.8078, 46.53802,
    45.08905,
  105.1592, 106.0084, 105.0161, 101.6408, 98.80224, 97.22235, 96.42387,
    95.73626, 91.93635, 93.3325, 94.14024, 93.10714, 93.68208, 93.06824,
    85.461, 74.15163, 71.00104, 75.56379, 77.67391, 73.73681, 68.99277,
    64.17552, 58.50844, 52.28091, 48.78102, 47.68568, 46.33887, 45.71909,
    45.47595, 44.77143,
  99.53284, 96.42339, 94.23776, 91.45171, 91.4055, 95.07713, 97.10199,
    96.51611, 92.55217, 92.26212, 89.26173, 84.77995, 84.69221, 86.7523,
    86.14647, 83.729, 78.71364, 75.33154, 73.58816, 68.81007, 59.52983,
    56.32335, 50.30428, 47.36223, 47.23267, 46.86985, 45.92978, 44.9836,
    44.44144, 44.0733,
  87.4753, 88.1162, 88.45341, 87.3701, 85.92851, 86.66524, 87.67916,
    83.90823, 79.18842, 75.56612, 74.52374, 72.0288, 71.52367, 74.7686,
    72.81859, 71.51019, 70.44202, 65.43649, 62.28008, 57.87144, 52.20504,
    51.39563, 47.83824, 46.8691, 47.07836, 46.89247, 45.95235, 45.06393,
    44.40329, 43.99876,
  77.32034, 75.57872, 74.51621, 73.97754, 73.40827, 72.71465, 72.74507,
    73.28793, 71.56947, 68.79768, 65.73456, 68.85994, 72.97595, 70.83096,
    66.88164, 64.21683, 61.26753, 59.154, 58.77522, 56.74341, 51.52458,
    51.17157, 48.17774, 47.00783, 47.031, 46.99022, 45.69495, 44.52217,
    44.1698, 43.95438,
  66.11815, 66.07078, 65.12368, 65.83534, 66.28156, 67.14819, 67.9946,
    69.36163, 70.14351, 68.85413, 71.48724, 74.68474, 74.20594, 73.02341,
    68.57274, 64.33266, 59.84779, 58.88527, 59.79132, 56.88491, 51.44133,
    50.48476, 48.58386, 47.71854, 46.81892, 46.13223, 45.28196, 44.09108,
    43.91597, 43.77751,
  72.8948, 69.29325, 63.60958, 60.83197, 62.22745, 62.3623, 63.2095,
    64.30773, 64.38638, 65.57812, 68.42094, 67.34192, 62.75832, 63.36092,
    62.23683, 63.01513, 67.02996, 70.77066, 70.0734, 64.8757, 56.72674,
    51.8338, 49.21964, 48.16769, 46.8227, 45.81732, 45.07566, 44.11093,
    43.84763, 43.75532,
  72.84441, 67.89205, 61.46579, 57.5933, 58.35916, 58.46052, 59.10973,
    60.06935, 61.79973, 64.80576, 65.52679, 62.03562, 61.83104, 61.53733,
    60.89135, 61.46833, 64.50459, 68.19006, 68.03548, 64.95623, 59.58265,
    54.21363, 50.53174, 49.34749, 47.95531, 46.27301, 45.25668, 44.3401,
    43.85249, 43.77873,
  69.64397, 65.47341, 59.11159, 55.76553, 56.43428, 56.75837, 57.5857,
    58.90916, 60.99682, 63.13725, 61.90148, 59.56446, 61.6574, 61.50768,
    60.22368, 59.3792, 59.7664, 60.19322, 59.98022, 58.18588, 56.51676,
    55.81058, 53.61856, 51.29861, 49.04186, 46.80498, 45.28704, 44.3541,
    43.83746, 43.77755,
  67.30287, 64.31326, 58.57854, 56.21749, 57.06474, 56.79306, 57.95053,
    58.98537, 61.16647, 61.84125, 58.77753, 56.84552, 57.88742, 57.42377,
    56.45191, 56.04799, 55.89346, 55.91057, 56.018, 55.62056, 55.09755,
    54.87239, 54.76166, 52.97005, 50.09174, 47.17511, 45.60117, 44.66208,
    43.91037, 43.76479,
  66.24078, 64.83658, 58.73374, 56.72113, 58.84672, 59.43869, 59.13818,
    57.73871, 57.88847, 56.76154, 53.52677, 53.5305, 54.1525, 54.51934,
    54.27885, 54.99393, 55.54498, 54.93147, 54.3667, 53.73249, 53.19115,
    52.84632, 52.25328, 51.52555, 51.17685, 48.71256, 46.48827, 45.60717,
    44.55384, 43.86127,
  68.71098, 68.71532, 64.33774, 62.46895, 62.86597, 62.0609, 62.02303,
    61.39463, 62.4455, 60.12562, 57.51974, 58.91228, 60.14214, 61.0732,
    60.79509, 60.82382, 60.57678, 58.71963, 55.94903, 54.23865, 53.32278,
    53.14252, 52.13094, 51.1292, 51.78195, 52.01701, 49.70478, 46.67861,
    45.54811, 44.34678,
  71.78951, 70.11309, 63.68787, 60.72713, 60.72266, 60.20774, 61.1062,
    63.64475, 66.95283, 64.3942, 61.4537, 63.75175, 65.36106, 65.87591,
    65.03293, 64.4649, 63.24532, 61.47071, 59.14587, 57.18441, 56.01703,
    54.89683, 52.90849, 51.70118, 52.52538, 53.69683, 52.95187, 49.43782,
    47.24147, 45.47821,
  75.10088, 74.77441, 67.80971, 62.63015, 61.67191, 61.70737, 64.74789,
    68.80652, 69.26174, 65.7393, 65.31291, 67.25074, 68.80935, 67.687,
    65.61168, 64.9464, 63.92021, 62.58778, 60.96328, 59.17958, 58.02135,
    56.4901, 53.81448, 52.52584, 53.10452, 53.22475, 53.17827, 50.46429,
    46.59569, 45.07169,
  76.49014, 74.90211, 68.61683, 64.13643, 63.30342, 62.48678, 65.83885,
    67.79079, 66.70557, 65.00305, 66.28333, 68.01516, 68.92284, 67.6105,
    65.74493, 64.8959, 63.81322, 62.81973, 61.58545, 60.79777, 60.87592,
    61.0182, 59.53911, 57.72289, 57.15255, 56.58637, 56.2977, 53.44843,
    47.15251, 44.23558,
  75.62444, 74.35561, 70.4012, 69.08309, 69.66801, 68.87825, 68.79878,
    67.56974, 64.78014, 64.98462, 66.05074, 67.96444, 69.3518, 68.96059,
    68.26522, 67.30255, 66.0864, 65.75842, 65.91185, 65.69003, 64.31471,
    62.27657, 59.54151, 58.16289, 58.01156, 57.58248, 56.76926, 56.0487,
    52.05473, 45.58302,
  68.17369, 68.32964, 68.73515, 69.40958, 71.56056, 73.13876, 70.22675,
    65.0444, 62.98649, 63.19139, 62.85012, 63.56551, 64.87444, 66.1442,
    67.01072, 66.63486, 65.25547, 64.02522, 61.83911, 59.26992, 57.95159,
    56.62172, 54.8748, 53.79971, 54.02964, 54.33683, 53.32587, 51.10125,
    49.40124, 46.51815,
  64.03675, 64.71331, 64.80099, 64.63045, 67.00668, 71.00488, 71.1785,
    65.22581, 62.27896, 63.27598, 63.7584, 64.72664, 65.01566, 64.32375,
    63.12998, 61.27227, 57.86614, 55.14979, 53.86102, 52.32255, 51.10221,
    51.01018, 50.83764, 50.34514, 50.31842, 50.58533, 49.6655, 47.53285,
    45.76063, 44.09959,
  50.66149, 50.63673, 50.72895, 50.75591, 50.68582, 50.7068, 50.81607,
    51.04655, 51.27661, 51.5408, 52.22111, 52.24965, 51.15467, 51.25727,
    51.23361, 50.95073, 51.01164, 51.1632, 51.42285, 52.00277, 52.17879,
    51.42529, 51.53946, 52.85882, 54.48558, 54.8163, 55.89914, 57.31615,
    53.13029, 51.36053,
  51.50708, 51.51947, 51.35657, 51.64883, 51.40302, 51.3292, 51.61941,
    51.98881, 52.3095, 52.6734, 53.14803, 53.50389, 53.40283, 52.52364,
    51.95064, 52.08256, 51.59571, 51.85223, 52.32216, 52.61347, 52.3662,
    52.42896, 54.53825, 59.67484, 64.3266, 60.73076, 55.55414, 58.31747,
    53.95823, 51.97265,
  51.41901, 51.30239, 51.30193, 51.32259, 51.26232, 51.35476, 51.56709,
    51.78136, 51.99955, 52.23917, 52.52591, 52.88981, 53.0266, 53.10197,
    53.05511, 52.28032, 52.58856, 53.68859, 54.82735, 57.39853, 62.61359,
    70.06334, 74.28507, 74.23077, 72.5871, 66.90988, 62.43211, 58.0001,
    54.02332, 52.52107,
  50.95698, 50.92195, 51.49678, 52.03012, 52.4529, 53.08835, 53.23079,
    53.26087, 53.64529, 54.09466, 54.33327, 54.73335, 54.61095, 54.28553,
    55.56242, 56.85143, 57.40396, 58.98895, 63.53575, 69.94005, 78.53739,
    80.84587, 76.18938, 75.83753, 71.35969, 69.24794, 67.62582, 59.83841,
    53.30706, 51.44828,
  51.46209, 51.38519, 52.50494, 53.49232, 54.12936, 54.42112, 54.54092,
    54.28395, 54.15316, 53.55241, 52.404, 52.21884, 52.74512, 54.26806,
    56.69901, 60.12296, 62.87153, 65.7336, 71.66511, 78.54012, 79.15047,
    70.61967, 66.73761, 69.13792, 69.87063, 69.13231, 68.36464, 73.51992,
    71.62365, 58.28121,
  51.75019, 52.42773, 53.59505, 54.24301, 53.02055, 51.64412, 51.29281,
    51.00599, 51.76201, 54.20156, 59.03192, 69.27726, 79.27574, 79.80606,
    83.46358, 87.282, 88.32045, 87.42899, 83.95201, 80.68565, 71.66246,
    62.67097, 66.28614, 69.74617, 73.42379, 74.60548, 76.17626, 86.31038,
    82.05216, 56.86142,
  51.09066, 51.67157, 52.87559, 54.13736, 55.05998, 58.68338, 68.00751,
    79.43443, 84.84232, 86.56378, 90.06946, 88.98203, 84.12097, 85.31226,
    86.54935, 87.17654, 86.99449, 82.12982, 76.07891, 72.53139, 67.70406,
    66.60845, 70.92102, 74.86582, 76.7011, 75.96246, 79.63503, 84.94669,
    71.94527, 50.50704,
  52.60463, 55.58272, 60.17421, 66.06524, 72.30847, 84.25158, 93.38141,
    88.81273, 83.9096, 84.16795, 81.07021, 76.06351, 72.4926, 71.96155,
    71.45348, 71.80627, 71.78622, 69.87148, 67.80997, 68.05082, 68.51141,
    70.24129, 73.37414, 75.75389, 75.26493, 76.39906, 81.65264, 79.49024,
    63.63084, 50.43486,
  62.47385, 68.29863, 74.17787, 80.00467, 87.06538, 90.98743, 82.19418,
    75.57578, 74.09146, 71.84646, 69.21381, 67.50967, 67.973, 70.9857,
    72.34379, 68.76383, 70.00241, 72.72383, 73.53738, 72.34869, 72.01704,
    75.26493, 79.05071, 78.79953, 77.76088, 83.23602, 85.2311, 72.94446,
    53.3754, 51.02126,
  78.11652, 84.94804, 84.03899, 86.21481, 88.73745, 82.36192, 65.46944,
    67.75658, 67.10242, 68.9738, 72.11815, 75.46091, 75.80503, 75.48283,
    74.51985, 76.4361, 79.2491, 80.51237, 79.93225, 80.16708, 81.06973,
    80.03982, 77.93029, 74.80426, 79.10672, 87.20397, 80.83978, 60.1073,
    50.61916, 50.6247,
  82.64323, 85.23656, 84.51871, 82.05991, 83.8829, 75.43182, 67.81336,
    73.28999, 77.59072, 80.25336, 76.25546, 69.23641, 68.18786, 68.89056,
    69.83934, 72.02705, 74.02782, 74.81782, 75.6273, 78.07061, 81.60822,
    79.03677, 72.998, 72.37331, 78.86235, 78.41471, 62.75824, 51.11538,
    51.4775, 50.50001,
  83.89033, 75.99545, 80.37798, 85.13988, 82.26237, 75.20224, 80.29491,
    76.53722, 71.85668, 71.86404, 67.41223, 64.39588, 66.90368, 67.78182,
    66.98222, 68.58518, 69.02504, 69.81262, 70.57057, 72.58301, 76.78045,
    76.5862, 73.07895, 78.70865, 81.0943, 67.80138, 51.53243, 52.90833,
    51.75272, 50.8438,
  94.61402, 96.92799, 100.8552, 103.0057, 103.3304, 101.3007, 87.39253,
    74.07153, 79.2828, 73.4664, 70.20435, 71.14213, 76.39561, 78.69603,
    74.32024, 66.13116, 67.95597, 69.10556, 70.06449, 72.55501, 76.771,
    78.27438, 76.37102, 72.68242, 68.38544, 60.25444, 52.35278, 54.0488,
    52.73969, 51.54064,
  100.4451, 104.4327, 105.7851, 103.5027, 100.5401, 97.2788, 94.6793,
    93.93141, 87.21329, 88.97705, 93.60603, 93.08605, 93.07297, 92.60117,
    85.77981, 75.74287, 74.75761, 80.86373, 84.58272, 81.15828, 78.01103,
    73.70117, 67.30501, 60.60053, 56.11188, 54.41938, 53.07096, 52.57179,
    52.17485, 51.47787,
  102.0296, 101.8484, 99.04683, 93.76183, 89.29721, 91.40133, 95.21243,
    95.26984, 92.39038, 93.5043, 91.76306, 87.38803, 86.90285, 88.78413,
    89.51135, 89.43034, 85.82419, 84.66698, 83.41676, 77.77059, 68.12992,
    64.0772, 57.52816, 53.9418, 53.91274, 53.71836, 52.84655, 51.83477,
    51.29099, 50.85938,
  95.31721, 91.37167, 89.09196, 87.42923, 87.71119, 90.04788, 91.91135,
    88.78711, 84.39851, 80.60945, 78.98567, 77.25378, 78.07936, 82.21545,
    81.59262, 80.68921, 79.62759, 74.68137, 70.55075, 65.05527, 59.19349,
    57.3828, 53.73086, 53.02817, 53.75323, 53.7987, 52.76904, 51.85317,
    51.20814, 50.77579,
  84.92871, 83.04456, 82.67818, 82.52029, 81.91135, 80.00682, 78.84469,
    78.57516, 76.42334, 73.85754, 71.8429, 74.79339, 78.73109, 77.31116,
    73.43446, 70.78014, 68.08512, 65.45302, 64.10491, 61.40152, 57.08234,
    56.68904, 54.01453, 53.12064, 53.62988, 53.84123, 52.57458, 51.44202,
    51.01595, 50.75939,
  76.76167, 76.68251, 75.18039, 74.27234, 72.82573, 72.05245, 72.0329,
    73.13988, 73.80962, 72.9501, 75.21667, 77.85324, 77.3056, 75.30073,
    71.052, 67.52076, 63.86563, 62.82109, 63.56691, 61.22391, 56.95961,
    56.45541, 54.62635, 53.84785, 53.41533, 52.9454, 52.11248, 51.01629,
    50.7193, 50.56998,
  81.13763, 77.18536, 70.62167, 66.90887, 67.53699, 67.57961, 68.52151,
    69.53847, 69.62956, 70.56673, 72.61336, 70.96527, 66.25768, 65.22021,
    63.24474, 63.47844, 67.07862, 71.06225, 71.59737, 67.93423, 61.97108,
    57.93188, 55.50749, 54.58003, 53.45405, 52.6482, 51.92544, 50.93504,
    50.59997, 50.52287,
  79.70915, 74.04466, 67.25999, 63.36505, 64.16138, 64.10461, 64.40744,
    64.56873, 64.98546, 66.54503, 66.40665, 62.9003, 61.98852, 61.39056,
    61.21188, 62.73797, 67.04939, 71.92291, 72.64248, 70.1916, 65.4369,
    60.04005, 56.4896, 55.59484, 54.4264, 53.06429, 52.06332, 51.07299,
    50.5871, 50.54759,
  75.72977, 71.12467, 64.26434, 60.33927, 60.32212, 59.81024, 59.71255,
    60.04318, 61.14847, 62.51476, 61.46292, 60.23239, 62.91913, 63.87513,
    64.04389, 64.81831, 66.48471, 67.65146, 67.09, 64.4325, 61.92588,
    60.57676, 58.75356, 57.02054, 55.43364, 53.68877, 52.18316, 51.14883,
    50.59902, 50.54433,
  72.12246, 68.53391, 61.66901, 58.05629, 57.95983, 57.09129, 57.91453,
    59.10946, 61.44159, 62.77986, 61.39687, 61.28454, 63.50856, 64.15059,
    63.90519, 63.65197, 63.27965, 62.89432, 62.27951, 61.14583, 60.38183,
    60.27847, 60.24843, 58.69694, 56.40387, 54.00159, 52.60203, 51.56509,
    50.6914, 50.52826,
  69.46436, 66.57075, 59.75298, 57.2706, 58.99049, 59.70145, 60.21901,
    60.27776, 61.49877, 61.37743, 59.5078, 60.10535, 60.97782, 61.11659,
    60.62805, 60.90263, 61.23454, 60.84855, 60.38275, 59.91932, 59.6078,
    59.37293, 58.6949, 57.54535, 56.93919, 54.87613, 53.14214, 52.36622,
    51.26748, 50.6095,
  69.93893, 68.879, 64.13719, 62.75109, 63.63913, 63.34578, 63.90734,
    64.08471, 65.27107, 63.59044, 61.66521, 63.08165, 64.29613, 64.75758,
    64.48876, 65.0941, 65.28525, 64.08482, 62.09009, 60.65839, 59.80383,
    59.46836, 58.27866, 56.93582, 57.18065, 57.21861, 55.61926, 53.34798,
    52.18157, 51.0716,
  73.68118, 71.90224, 65.22156, 62.54541, 62.35465, 61.96552, 63.00741,
    65.36008, 68.20558, 66.16257, 63.91519, 66.36058, 68.5782, 69.29573,
    68.95087, 69.18478, 68.29809, 66.96091, 65.05004, 63.36356, 62.08272,
    60.66972, 58.68046, 57.32004, 57.86929, 58.79267, 58.33859, 55.59394,
    53.6909, 52.02042,
  75.13229, 74.11383, 67.2507, 62.66808, 61.81004, 61.92126, 64.58964,
    68.62431, 69.92934, 67.34227, 67.33076, 69.78067, 71.95736, 71.62621,
    70.14668, 69.89352, 69.27603, 68.13615, 66.75349, 65.29394, 63.83218,
    61.97562, 59.48293, 58.23043, 58.66999, 58.7245, 58.69014, 56.41845,
    53.29464, 51.76232,
  74.9377, 72.98625, 67.05925, 63.26725, 62.89392, 62.54086, 65.73782,
    68.27005, 68.34055, 67.43844, 69.0151, 71.08826, 72.42106, 71.29343,
    69.79688, 69.5809, 68.99759, 67.9996, 66.69235, 65.70531, 65.36548,
    65.04732, 63.43105, 61.70408, 61.21925, 60.92681, 61.04571, 58.77992,
    53.52198, 51.01633,
  73.61161, 72.01114, 68.16253, 66.94305, 67.98283, 68.0724, 68.78933,
    68.55724, 67.06422, 67.63406, 69.0977, 70.99174, 72.37757, 72.03416,
    71.23978, 70.6731, 70.05748, 69.55966, 69.53731, 69.57431, 68.51196,
    66.71377, 64.07959, 62.64569, 62.43645, 62.08194, 61.66294, 60.91704,
    57.32598, 51.98739,
  67.20854, 67.50814, 67.86879, 68.64656, 71.04755, 72.80032, 70.75327,
    66.75755, 65.374, 65.73264, 65.752, 66.53529, 67.85824, 69.34846,
    70.4031, 70.72685, 70.41388, 69.85336, 68.3756, 66.44467, 65.02652,
    63.57893, 61.775, 60.76202, 60.73618, 60.47133, 59.51356, 57.70016,
    56.049, 52.98806,
  64.14185, 64.70633, 65.13198, 65.41983, 67.63107, 71.21944, 71.51385,
    66.76452, 64.63237, 65.65778, 66.26292, 67.1992, 67.89598, 68.26924,
    68.22395, 67.38528, 65.07579, 63.24395, 62.20229, 60.49656, 59.14922,
    58.85303, 58.49181, 57.99701, 57.5162, 57.04013, 56.02665, 54.46105,
    52.9208, 51.07145,
  5.686986, 4.910253, 5.251091, 5.404831, 5.501674, 5.619334, 5.860106,
    6.194597, 6.715848, 7.699177, 9.506939, 11.59907, 13.00764, 16.13237,
    19.86292, 24.04504, 28.89959, 34.70696, 39.23046, 44.09304, 48.94336,
    52.90406, 55.77557, 57.65443, 57.74449, 55.16594, 53.41701, 56.20493,
    49.90709, 47.20975,
  5.020844, 4.506449, 4.661834, 5.223485, 5.469644, 5.625019, 5.992643,
    6.247455, 6.569919, 7.241548, 8.715463, 11.2284, 14.35097, 16.86487,
    20.14829, 25.24465, 30.6743, 35.13398, 39.97707, 45.31134, 50.04124,
    54.12032, 57.04714, 58.86016, 59.56696, 58.94511, 52.88607, 54.46078,
    50.09934, 47.87818,
  7.746788, 7.748677, 8.629617, 9.216511, 9.996878, 10.88639, 11.64337,
    12.31546, 12.7569, 13.02222, 13.46245, 14.52762, 16.33568, 18.8884,
    21.94329, 24.83655, 30.07729, 36.01698, 41.13844, 46.69144, 51.97435,
    56.28952, 59.19677, 60.47001, 60.46811, 59.87526, 59.36316, 55.75022,
    49.15464, 47.95337,
  10.71044, 11.26772, 12.63687, 13.70317, 14.42826, 14.92995, 15.06426,
    15.19388, 15.5129, 16.12653, 17.16567, 18.48507, 20.16817, 22.5421,
    25.48313, 28.66501, 32.28275, 36.21929, 41.25709, 46.87196, 52.33575,
    56.59329, 58.95657, 60.66638, 60.79853, 60.78025, 60.75185, 59.59021,
    57.59415, 48.60072,
  13.40433, 14.29502, 15.17237, 15.14778, 15.20231, 15.20075, 15.25733,
    15.3171, 15.64508, 16.42946, 17.71356, 19.51921, 21.56079, 23.96846,
    26.78772, 29.96055, 33.54876, 37.62993, 42.43695, 48.00347, 52.7635,
    56.03566, 58.67632, 60.18731, 60.61752, 60.56139, 60.34118, 61.12523,
    60.68764, 58.63219,
  12.89332, 14.54023, 15.41841, 15.63369, 15.75024, 15.76469, 15.98173,
    16.11867, 16.16278, 16.54673, 17.60788, 19.41185, 22.03968, 24.65789,
    27.6482, 31.08888, 35.22501, 39.46636, 43.9493, 49.15202, 53.38553,
    56.03246, 59.01812, 60.16843, 60.39432, 60.07722, 59.52233, 60.12252,
    60.06732, 52.10377,
  13.20255, 14.13465, 15.40569, 15.6283, 15.91053, 16.18099, 16.58376,
    17.06345, 17.42595, 17.74923, 18.46547, 19.42393, 18.92577, 22.57845,
    26.39174, 30.02615, 34.08821, 38.84033, 43.51084, 48.96241, 53.5572,
    57.01382, 59.31102, 60.48641, 60.51318, 59.80912, 59.6361, 59.76904,
    59.07281, 45.55799,
  16.34116, 15.38822, 15.82288, 15.89583, 16.0324, 16.47622, 16.81963,
    15.87257, 13.29423, 16.54425, 17.64405, 18.69378, 20.93681, 23.83142,
    26.8852, 30.18889, 34.3839, 39.15465, 44.01506, 49.06743, 53.74297,
    57.32275, 59.64122, 60.62209, 60.32662, 59.98911, 60.13287, 59.73306,
    58.3495, 45.86708,
  19.31394, 17.58898, 17.34515, 17.03749, 16.81419, 16.72268, 15.75105,
    14.82291, 15.17178, 15.82318, 17.86666, 19.7563, 21.83151, 24.63745,
    27.87386, 30.57068, 34.5912, 39.92225, 45.22454, 50.02819, 54.42692,
    57.92799, 59.91667, 60.3574, 60.05904, 60.34573, 60.15995, 59.13625,
    46.19075, 46.50605,
  24.35308, 22.34584, 20.87052, 19.75785, 19.18671, 18.19762, 16.38756,
    16.63682, 16.55854, 17.04225, 18.27353, 20.53269, 22.79886, 24.77364,
    27.16698, 30.83505, 35.05499, 39.78656, 44.94453, 50.3588, 55.34849,
    58.45787, 59.42526, 59.151, 59.52908, 59.9388, 59.5248, 53.16975,
    45.81164, 45.48313,
  29.06946, 26.59424, 26.56193, 24.23845, 23.03114, 21.1766, 19.56744,
    18.57541, 18.3452, 18.9579, 19.52754, 20.77706, 22.41515, 24.74231,
    27.46906, 30.77222, 34.69046, 39.17672, 44.11744, 49.35411, 55.01583,
    58.30055, 59.07933, 59.11308, 59.50309, 59.17788, 55.22983, 46.37525,
    46.82429, 45.60633,
  29.56041, 27.63542, 30.20484, 30.53012, 29.20329, 25.47645, 22.20302,
    19.17261, 17.98212, 18.54716, 19.6266, 21.20762, 23.67381, 25.73769,
    28.11849, 31.60259, 34.95578, 39.35329, 44.23277, 49.14533, 54.03377,
    57.82557, 58.77134, 59.50041, 59.79539, 58.85428, 46.47094, 51.17453,
    47.53078, 46.33633,
  19.98142, 21.43791, 23.79935, 26.74713, 28.81831, 28.30963, 21.96919,
    16.7093, 20.3556, 19.14936, 20.60518, 21.68966, 23.8395, 26.19635,
    28.81439, 31.16315, 35.23702, 39.71585, 44.59948, 49.562, 54.08524,
    57.12297, 58.44295, 56.94277, 56.65717, 55.45094, 47.46046, 49.10436,
    48.58488, 47.2107,
  15.98352, 14.90657, 15.08722, 15.35816, 15.90584, 16.58791, 17.46261,
    18.79219, 17.78392, 18.9727, 20.72811, 22.69567, 24.52234, 26.48684,
    29.22211, 31.86354, 34.89312, 40.20463, 45.52378, 50.25662, 53.87724,
    56.53804, 55.0801, 50.15079, 47.04612, 47.26972, 46.76472, 46.33673,
    46.56311, 46.59161,
  16.8762, 12.65333, 16.10653, 16.36876, 16.6439, 16.79065, 17.10779,
    17.30961, 17.7799, 19.04753, 20.69917, 22.5964, 24.7012, 27.04826,
    29.0518, 31.69377, 35.48128, 38.88239, 44.49389, 49.84079, 50.29194,
    52.9351, 50.60431, 48.39657, 48.70442, 47.79458, 47.07204, 46.51464,
    45.96682, 45.78548,
  10.85111, 12.11484, 13.8974, 15.9558, 16.39607, 16.96313, 17.62928,
    17.93121, 18.47812, 20.06941, 22.36614, 24.26666, 26.12291, 27.79859,
    29.8364, 32.42488, 35.28074, 38.90912, 41.28643, 45.22426, 45.77689,
    49.08521, 48.85764, 48.58686, 48.51107, 47.83424, 47.01117, 46.59083,
    46.06937, 45.82538,
  7.884311, 6.440423, 8.012371, 9.724138, 11.68037, 14.19202, 16.36194,
    17.10804, 18.27553, 20.06986, 22.15384, 24.94566, 28.10516, 30.06624,
    32.1439, 34.37522, 36.87567, 40.52875, 43.88256, 46.52112, 46.05558,
    49.20633, 49.10973, 48.66258, 48.47641, 48.01865, 46.9567, 45.95828,
    45.71695, 45.6953,
  10.93333, 7.989293, 6.91992, 7.390333, 8.688113, 9.925195, 11.37214,
    12.94439, 15.42585, 17.85376, 20.52269, 23.60975, 26.5384, 30.58555,
    33.95603, 36.53492, 39.31649, 43.56584, 48.70446, 52.739, 49.36916,
    49.57482, 49.24908, 48.99936, 48.29884, 47.76753, 47.03799, 45.83325,
    45.52168, 45.52676,
  24.79983, 17.17862, 9.895409, 4.698983, 6.758984, 6.899568, 7.921725,
    9.061921, 10.26614, 12.44866, 15.82289, 18.36707, 20.18737, 26.10368,
    32.0377, 36.05449, 40.56902, 46.22243, 52.17437, 56.52546, 58.24443,
    53.69049, 50.77672, 50.48745, 49.04778, 48.1957, 47.31833, 46.06786,
    45.50235, 45.56718,
  24.68853, 17.92932, 10.34395, 5.132272, 6.623139, 6.847507, 7.825748,
    8.997497, 10.86353, 13.78374, 15.94872, 15.68005, 18.36129, 20.61179,
    24.07048, 28.70472, 35.31672, 43.33624, 49.87867, 54.74022, 58.08796,
    56.87991, 53.18009, 52.00756, 50.37659, 48.78678, 47.62227, 46.23359,
    45.47036, 45.57898,
  27.0265, 20.6126, 12.793, 7.523089, 8.454763, 8.295538, 9.026941, 10.03205,
    11.7878, 13.76138, 14.4251, 15.07934, 19.0846, 21.68739, 24.29864,
    27.99921, 33.18184, 39.41841, 45.62543, 50.52138, 54.32111, 56.71784,
    55.78598, 53.81404, 51.74495, 49.51364, 47.77795, 46.27225, 45.47566,
    45.58668,
  27.66155, 23.94781, 16.72484, 12.48349, 13.9924, 13.28568, 13.83472,
    14.15036, 15.76434, 16.96113, 16.47488, 17.49532, 20.64098, 23.46364,
    26.21127, 29.87347, 34.22711, 39.37983, 44.71846, 49.00635, 52.52484,
    54.65541, 56.01203, 55.81826, 53.84196, 50.55791, 48.37925, 46.90551,
    45.67321, 45.56276,
  28.02806, 24.9525, 19.96999, 16.66092, 19.47563, 20.4119, 21.05463,
    20.79356, 21.51736, 22.08477, 22.21966, 24.92826, 27.7824, 30.38103,
    32.56233, 35.80354, 39.62344, 43.16834, 47.10943, 50.44974, 53.00163,
    54.50359, 55.09758, 55.51065, 55.89699, 53.01901, 49.79326, 47.98592,
    46.60461, 45.74993,
  28.24172, 24.90917, 21.53369, 19.62416, 21.0969, 21.73333, 23.07538,
    24.6354, 26.47417, 27.66581, 28.45055, 32.57153, 36.22071, 39.21879,
    41.46067, 44.37531, 47.71777, 50.37983, 52.88197, 55.38419, 56.98788,
    57.11427, 56.39562, 55.99693, 56.60181, 56.23927, 53.48376, 49.54326,
    47.96143, 46.6142,
  28.21872, 23.86323, 19.58009, 16.26617, 18.37068, 19.48039, 21.45997,
    23.53158, 25.64062, 26.94255, 27.72034, 31.96036, 35.94642, 39.2734,
    41.56025, 44.63697, 47.9743, 51.77107, 55.2805, 57.99051, 59.56151,
    59.46487, 57.56727, 55.92542, 56.08381, 55.93426, 54.98316, 51.26845,
    48.74303, 47.50411,
  29.74883, 25.70071, 21.98991, 18.423, 18.94463, 19.61478, 22.32447,
    24.51343, 26.30583, 27.13646, 29.58696, 32.8994, 36.60406, 39.55091,
    41.71615, 44.73687, 48.10226, 51.43841, 55.2756, 58.95031, 61.36089,
    61.97703, 60.18505, 58.06019, 57.64602, 56.52936, 55.52646, 52.42204,
    48.12961, 46.90124,
  36.66796, 33.02876, 29.45851, 26.19407, 26.43933, 25.59901, 27.63623,
    29.15738, 29.74039, 30.83238, 34.04524, 37.86547, 41.46089, 43.92442,
    45.11266, 46.97885, 48.9929, 51.59935, 54.64661, 58.10196, 60.77976,
    62.2373, 61.65368, 60.1389, 59.68252, 58.90977, 58.50812, 56.04008,
    49.91084, 46.45994,
  47.36049, 45.60385, 42.53902, 41.01682, 41.93517, 42.17682, 41.15185,
    40.29282, 39.36597, 40.1735, 41.48283, 43.79621, 46.83624, 49.01,
    49.66259, 50.60099, 51.14784, 52.19516, 54.41383, 57.08583, 57.96077,
    57.85931, 56.69515, 55.85422, 56.20671, 56.12938, 55.89647, 55.61549,
    53.16755, 47.98925,
  48.62642, 49.58234, 51.62217, 52.4432, 53.33804, 54.37411, 53.74615,
    49.23578, 47.79808, 48.2155, 47.8783, 48.0424, 48.54724, 49.26962,
    49.65778, 49.91533, 49.66806, 49.76172, 50.03124, 50.29787, 51.00749,
    52.00948, 52.20329, 51.51639, 51.68641, 51.80852, 51.29696, 49.83971,
    49.22277, 48.1018,
  50.30959, 50.97044, 51.51668, 51.54282, 52.77133, 55.47184, 55.82205,
    52.09609, 49.66093, 50.58484, 51.09021, 51.44766, 51.54216, 51.20771,
    50.66577, 50.07973, 48.91417, 47.53513, 47.47819, 47.44534, 47.12215,
    47.86505, 48.72958, 49.15038, 49.05399, 49.31833, 49.13646, 47.91067,
    46.69058, 45.78838,
  26.94531, 28.79697, 31.14576, 33.49156, 35.88435, 38.43791, 40.91066,
    43.59188, 46.48146, 49.38498, 52.21947, 54.75325, 56.56475, 58.07412,
    59.11459, 59.80459, 60.19386, 60.55485, 60.88198, 61.25385, 61.61562,
    61.82612, 62.05019, 62.32216, 62.27929, 61.72904, 55.1618, 58.43084,
    53.9279, 50.67608,
  25.9926, 27.73534, 30.2722, 33.00135, 35.68222, 38.55476, 41.38116,
    44.32292, 47.19474, 50.05813, 52.87903, 55.48951, 57.60751, 58.93471,
    59.67496, 60.12055, 60.33881, 60.6688, 61.06721, 61.65102, 62.33215,
    62.9966, 63.50921, 63.90809, 64.02246, 63.08311, 61.51264, 56.47723,
    53.1736, 51.07729,
  27.04335, 28.45731, 30.8935, 33.43484, 35.91854, 38.84218, 41.85413,
    45.00425, 48.08382, 50.91908, 53.58422, 55.97345, 58.04658, 59.49843,
    60.33026, 60.54138, 60.56399, 60.76748, 61.08595, 61.49333, 62.37013,
    63.46254, 64.17628, 64.57776, 64.46129, 64.16969, 63.46412, 61.89334,
    53.46812, 50.68051,
  27.58622, 29.29651, 31.89132, 34.29213, 36.60976, 39.03284, 41.79911,
    44.92439, 48.15725, 51.31076, 54.13868, 56.58595, 58.66953, 59.99702,
    60.84938, 61.25204, 61.15595, 61.08807, 61.42784, 61.86177, 62.53114,
    63.00944, 62.92455, 63.85622, 63.94294, 64.24763, 64.53027, 63.76242,
    62.16622, 53.58532,
  28.20707, 30.12738, 32.65877, 35.37699, 37.68621, 39.9351, 42.17167,
    45.06842, 47.90409, 51.03352, 54.05359, 56.78257, 59.28131, 60.82108,
    61.62251, 62.03724, 61.99316, 61.72869, 61.83469, 62.30692, 62.5086,
    62.14754, 62.61213, 63.393, 63.77874, 63.7676, 63.85509, 64.88198,
    64.50632, 62.07116,
  29.11242, 30.69729, 33.25322, 35.89508, 38.57008, 40.81339, 43.05351,
    46.00863, 48.5589, 51.01291, 53.76488, 56.51733, 59.32199, 61.07899,
    62.13309, 62.64626, 62.64062, 62.39373, 61.99964, 62.1886, 62.13984,
    61.88414, 62.88841, 63.65364, 63.99426, 63.83316, 63.43737, 63.98378,
    63.81058, 55.70567,
  31.91455, 32.28613, 34.25533, 36.35061, 38.9416, 41.42067, 43.73453,
    46.66688, 49.45734, 51.8628, 54.21686, 56.09101, 57.24179, 59.14982,
    60.40786, 61.24415, 61.67828, 61.46305, 60.97756, 61.15949, 61.44791,
    61.95766, 62.85269, 63.80067, 64.14546, 63.87136, 63.79247, 63.63227,
    62.58841, 48.88357,
  37.12477, 36.30582, 36.91078, 38.08792, 39.89585, 42.51383, 44.93424,
    46.04301, 47.89243, 50.43942, 52.66885, 54.8721, 56.92419, 58.83421,
    60.22185, 61.09438, 61.83455, 62.13523, 61.86799, 61.54637, 61.58706,
    62.01394, 62.78975, 63.57907, 63.76272, 63.98354, 64.10723, 63.26493,
    61.55677, 49.22178,
  43.1806, 42.95726, 42.17362, 41.98915, 42.58823, 44.06668, 44.80236,
    46.74834, 49.21696, 51.41726, 53.40873, 55.30057, 56.88221, 58.5496,
    60.09259, 60.65682, 61.43926, 62.41619, 62.92261, 62.64066, 62.43087,
    62.45397, 62.71233, 62.86588, 63.05922, 63.84623, 63.97651, 62.63206,
    49.07296, 49.90677,
  46.01138, 48.71947, 49.02081, 48.12653, 47.22503, 46.85196, 46.50164,
    48.29527, 50.26073, 52.63776, 54.34698, 56.02025, 57.26824, 58.21833,
    58.90958, 59.95872, 60.72014, 61.44593, 62.15617, 62.43786, 62.95802,
    62.81976, 62.5732, 62.17661, 62.59531, 63.00853, 62.77488, 56.94189,
    49.49631, 48.99886,
  43.88956, 47.20419, 51.87309, 53.53902, 53.25368, 51.20863, 50.18206,
    50.49266, 51.52769, 54.02611, 55.52136, 56.2786, 57.31036, 58.11058,
    58.81046, 59.46218, 60.0345, 60.52539, 61.06252, 61.42118, 62.31575,
    62.41952, 62.00794, 62.47583, 63.26147, 62.73396, 60.42387, 51.08257,
    50.60946, 49.29916,
  39.77637, 40.22305, 47.54536, 53.45941, 57.94791, 56.39341, 53.14189,
    50.87422, 52.57753, 53.80197, 55.81078, 57.10305, 58.64918, 59.3502,
    59.5085, 59.68075, 60.31066, 60.75472, 61.02296, 61.16501, 61.8146,
    62.02936, 61.44311, 62.03964, 63.08981, 62.54949, 49.49688, 56.13223,
    51.90195, 50.23499,
  33.86526, 36.25643, 39.23716, 44.97805, 51.36125, 55.97614, 53.41364,
    49.65201, 55.22406, 55.49118, 57.4817, 58.58071, 59.9959, 61.00226,
    61.15597, 59.87241, 60.47432, 61.25599, 61.56985, 61.35169, 61.78111,
    61.84105, 61.43388, 59.61056, 58.11706, 60.22854, 50.43747, 52.0004,
    52.44268, 51.10798,
  32.48954, 34.03394, 35.69549, 37.97969, 40.50003, 43.49757, 47.83146,
    52.46043, 53.44786, 56.05959, 58.38163, 60.25347, 61.24206, 62.04092,
    62.13877, 61.21836, 60.54539, 61.17014, 61.94487, 61.57573, 61.21653,
    61.18075, 59.87025, 54.09933, 49.89989, 50.28761, 50.36565, 49.48812,
    49.73775, 50.08976,
  30.86405, 28.82744, 34.94086, 38.10718, 40.86625, 43.79632, 46.39721,
    49.4127, 53.04777, 55.91563, 58.06374, 59.80432, 61.4284, 62.70251,
    62.88229, 62.78831, 61.77808, 60.76075, 60.56147, 60.69023, 57.54788,
    58.15745, 54.44763, 51.40746, 52.23162, 51.20301, 50.67115, 50.13251,
    49.41258, 49.22082,
  25.09248, 27.37398, 30.01168, 33.92278, 38.31995, 41.79883, 44.78892,
    47.84325, 51.04411, 54.50978, 57.34644, 59.54993, 61.41655, 63.1179,
    63.7211, 63.55879, 63.25869, 62.05835, 60.07006, 56.93894, 53.72594,
    54.22363, 52.60218, 51.68138, 51.60505, 51.13123, 50.32909, 49.88287,
    49.51735, 49.3382,
  28.74907, 27.30522, 30.09127, 32.94443, 36.06822, 39.81499, 43.65425,
    46.97357, 49.73051, 52.79333, 55.56465, 58.49073, 61.1851, 62.76482,
    63.76461, 64.52224, 64.84545, 64.53401, 63.52768, 62.08673, 55.21012,
    54.15364, 52.86554, 52.11579, 51.96167, 51.59393, 50.38737, 49.38054,
    49.16541, 49.17544,
  39.70834, 34.44183, 32.98649, 34.25887, 37.94659, 40.71543, 43.98954,
    47.08009, 50.36502, 52.64158, 55.48347, 57.98288, 59.7423, 61.40759,
    62.52565, 63.69944, 64.90956, 65.93213, 66.32684, 65.2891, 62.29029, 56,
    53.49633, 53.10803, 52.15516, 51.76788, 50.74926, 49.35787, 49.09072,
    49.04511,
  50.29086, 45.88889, 40.8825, 35.27399, 39.9067, 42.00313, 45.22206,
    48.43391, 51.69763, 54.85393, 57.33585, 58.91262, 57.70171, 58.0148,
    58.76278, 61.12763, 63.30802, 65.12449, 66.2807, 66.78413, 65.70363,
    62.0622, 55.80957, 55.27794, 53.54472, 52.62496, 51.38797, 49.70913,
    49.03408, 49.08915,
  49.82583, 47.0403, 43.09906, 39.30902, 43.12041, 45.07927, 48.24407,
    51.47356, 54.95277, 57.48281, 59.4106, 60.64256, 61.9731, 61.55066,
    60.04988, 59.1819, 59.95038, 62.5211, 63.85252, 64.12926, 64.57886,
    64.12592, 59.13111, 57.19501, 55.42627, 53.55252, 51.9174, 49.91705,
    48.95749, 49.10696,
  51.40824, 48.53653, 44.75804, 43.21329, 46.71569, 48.86251, 51.97685,
    54.90186, 57.62515, 59.96569, 61.6048, 62.33356, 64.08612, 64.74728,
    64.222, 63.39192, 62.88049, 63.24498, 63.18325, 62.38437, 62.37971,
    62.83015, 61.55895, 59.35522, 57.366, 54.64152, 52.28981, 50.16689,
    48.99345, 49.11084,
  53.7793, 51.0947, 47.46817, 45.98945, 49.49924, 51.73453, 54.64384,
    57.46093, 60.35324, 62.9903, 64.91882, 66.37897, 67.35817, 67.67803,
    67.56083, 67.17833, 66.40862, 65.42192, 64.73502, 63.20505, 62.01935,
    61.35712, 61.70457, 60.74302, 59.21906, 55.9432, 53.10404, 51.15394,
    49.43955, 49.08108,
  59.06155, 56.26011, 52.25483, 50.37395, 53.56702, 55.77406, 58.55276,
    61.13512, 63.771, 66.10052, 68.30468, 70.63679, 72.20528, 72.49001,
    71.99871, 71.49032, 70.71332, 69.75748, 68.59797, 66.92305, 65.17948,
    63.16713, 62.05098, 61.23545, 61.36625, 58.37989, 54.65811, 52.25431,
    50.58296, 49.43007,
  65.827, 62.3, 57.90867, 55.85733, 57.97878, 59.3544, 61.77401, 64.61471,
    67.60519, 69.37897, 71.13412, 73.8205, 76.60242, 77.67294, 76.71701,
    76.31897, 75.29884, 74.05215, 72.65141, 71.59974, 70.54884, 67.64999,
    64.65255, 62.84243, 62.79739, 61.51101, 58.16253, 53.62144, 51.85349,
    50.43307,
  71.73, 67.27274, 62.08315, 58.93114, 60.45253, 60.99279, 62.66894,
    65.29705, 68.00844, 69.29882, 70.65713, 72.9204, 75.54324, 76.66589,
    75.58899, 75.30608, 74.82377, 74.04754, 73.04054, 72.41858, 71.67394,
    69.29166, 65.83014, 63.58652, 63.29744, 62.00465, 60.13352, 55.43443,
    52.14523, 51.11826,
  74.86024, 70.26872, 65.10719, 61.59731, 61.47466, 60.98899, 63.53288,
    65.47873, 67.26559, 67.68815, 69.32034, 71.79266, 74.47131, 75.25615,
    74.01331, 73.71785, 73.40704, 72.75771, 72.0921, 71.83689, 71.0482,
    69.47549, 66.47472, 64.12784, 64.06533, 62.96541, 61.42163, 57.35645,
    52.24625, 50.59206,
  74.56284, 71.017, 66.12029, 63.02602, 62.95253, 60.9808, 61.79771,
    63.25474, 63.16888, 62.69279, 64.31325, 67.80414, 71.53111, 72.96498,
    71.99728, 71.01662, 69.96925, 69.25183, 68.74752, 68.84127, 68.46724,
    67.34731, 65.0252, 63.10653, 63.16522, 62.77396, 62.51199, 60.36523,
    54.6702, 50.57704,
  70.1312, 68.20763, 65.03832, 62.91704, 63.74385, 63.50564, 61.9926,
    60.89711, 59.65058, 59.28294, 59.24842, 60.79882, 63.84889, 66.16864,
    65.72639, 64.94269, 63.37241, 62.07447, 62.12955, 63.27235, 63.31014,
    62.48801, 60.2705, 58.75245, 59.12766, 58.76415, 58.26614, 57.92775,
    56.17079, 51.86616,
  56.20597, 57.33159, 58.90055, 60.32924, 61.51155, 62.90622, 61.40853,
    57.38593, 55.68965, 56.0369, 55.48936, 55.19565, 55.43122, 56.27164,
    56.45672, 56.18575, 55.13097, 54.04028, 53.48704, 53.38918, 53.85265,
    55.01558, 55.62835, 54.98706, 55.18001, 55.27748, 54.5545, 52.83158,
    51.85021, 51.23228,
  53.29411, 53.69349, 54.08334, 54.11512, 54.63123, 56.62034, 57.57109,
    54.69582, 52.6326, 53.29193, 53.5604, 53.59369, 53.47578, 53.32412,
    53.22197, 52.99022, 51.87556, 50.65805, 50.40532, 50.31412, 50.01805,
    50.50989, 51.51274, 52.17233, 52.07, 52.26057, 52.23087, 51.24214,
    49.98586, 49.24297,
  56.89373, 58.20198, 59.22911, 60.15856, 60.71752, 61.16445, 61.53268,
    61.79637, 62.03565, 62.30164, 62.68771, 63.04842, 63.39116, 63.8509,
    64.36266, 65.01199, 65.77038, 66.70823, 67.88787, 69.28837, 70.69602,
    72.11201, 73.26939, 73.7541, 68.55812, 60.47008, 54.66678, 57.22429,
    54.05024, 51.77423,
  56.2725, 57.58893, 58.71507, 59.73245, 60.40092, 60.88949, 61.29346,
    61.70523, 62.03233, 62.29337, 62.63763, 63.02853, 63.46492, 63.91514,
    64.37067, 64.96236, 65.67404, 66.58752, 67.7702, 69.21627, 70.98597,
    72.87096, 74.37133, 75.36063, 75.4388, 74.03624, 58.16865, 55.00742,
    53.5117, 52.03168,
  56.5313, 57.74689, 58.79159, 59.76507, 60.50381, 61.0647, 61.46794,
    61.90078, 62.35587, 62.72834, 63.07552, 63.47917, 63.86135, 64.34232,
    64.9259, 65.51714, 66.17365, 67.00011, 67.90085, 69.1638, 70.94686,
    73.07607, 74.86932, 75.96707, 76.01429, 75.11606, 73.9915, 61.5519,
    53.38259, 51.86279,
  56.66806, 57.81945, 58.84257, 59.73954, 60.49508, 61.16066, 61.56453,
    61.89868, 62.31581, 62.73954, 63.3505, 64.03128, 64.5573, 64.9005,
    65.43277, 66.10069, 66.72008, 67.35767, 68.34151, 69.56525, 70.97501,
    72.2799, 71.4041, 74.9642, 75.38984, 75.58624, 75.17625, 74.37084,
    66.2936, 54.14819,
  56.99311, 58.01778, 59.02461, 59.88253, 60.53427, 61.19605, 61.79828,
    62.07768, 62.26492, 62.59515, 63.22923, 64.35806, 65.4302, 65.9213,
    66.46685, 67.02834, 67.48894, 67.9277, 68.77335, 70.04694, 70.99875,
    69.26878, 67.24721, 69.2532, 71.99969, 75.02901, 74.96301, 75.79272,
    75.66185, 64.96685,
  57.63768, 58.37622, 59.45464, 60.2243, 60.73102, 61.23901, 62.05079,
    62.67067, 62.81397, 62.82872, 63.18547, 64.19806, 65.60072, 66.39803,
    67.1509, 67.74901, 68.0247, 68.48775, 68.95632, 69.87536, 70.62671,
    66.45596, 71.92462, 72.35598, 72.43903, 72.35114, 73.49461, 74.82111,
    74.92567, 57.17265,
  59.69137, 59.42025, 60.22397, 60.76582, 61.19458, 61.63029, 62.33084,
    62.75506, 63.13913, 63.24317, 63.48516, 63.6332, 63.55686, 64.55293,
    65.40559, 66.19341, 66.70076, 67.21453, 67.85656, 68.92545, 70.06824,
    69.13174, 72.11015, 74.67519, 75.05431, 74.8529, 74.80445, 74.66628,
    73.83667, 50.60371,
  64.04916, 62.29446, 62.02169, 61.92636, 62.03624, 62.52125, 62.8762,
    61.80593, 61.19708, 61.51334, 61.88489, 62.49633, 63.30774, 64.28323,
    65.17133, 65.91257, 66.79315, 67.64402, 68.30533, 69.09389, 69.55346,
    70.53272, 72.51588, 74.54548, 75.02242, 75.29404, 75.21372, 74.30595,
    65.08111, 50.8703,
  69.85909, 68.19962, 66.10807, 64.69744, 63.76001, 63.34581, 62.2281,
    62.24146, 62.23413, 62.06349, 62.24346, 62.66111, 63.16134, 64.11871,
    65.18917, 65.79623, 66.82148, 68.15532, 69.26039, 69.92693, 70.85083,
    71.88043, 72.92272, 73.68885, 74.44283, 75.26205, 75.30501, 74.04456,
    50.74389, 51.48063,
  72.90852, 74.1553, 72.51633, 70.20177, 67.73714, 65.38645, 63.19919,
    63.25544, 63.22138, 63.30623, 63.07491, 63.19523, 63.4473, 63.89449,
    63.66175, 63.44152, 63.92239, 65.55476, 67.81511, 69.94258, 71.25635,
    72.15223, 72.65906, 73.07803, 73.9978, 74.50014, 74.15562, 58.09682,
    50.91134, 50.91099,
  70.49814, 73.25034, 76.49734, 76.11615, 73.93314, 69.54546, 66.46061,
    64.75605, 64.02518, 64.71899, 64.17697, 63.55745, 63.62024, 64.01463,
    63.97973, 63.68427, 62.34233, 61.42056, 62.01423, 64.08218, 67.72567,
    69.57467, 71.73125, 73.42037, 74.72904, 74.5546, 61.55817, 52.07712,
    52.20882, 51.09561,
  66.08504, 66.21797, 71.82381, 75.97919, 77.44793, 74.05424, 69.31104,
    65.75684, 64.92337, 64.78786, 64.59533, 64.2921, 64.81149, 64.9661,
    64.86147, 65.39962, 66.41636, 66.23669, 63.76412, 62.88649, 65.39828,
    66.63451, 66.19422, 71.3557, 74.3499, 74.08759, 51.3167, 57.30709,
    53.11418, 51.8108,
  60.19374, 61.73723, 63.46363, 66.90176, 70.70201, 72.59879, 68.17089,
    64.5536, 67.19904, 66.18655, 66.03772, 65.51385, 65.98056, 66.36419,
    66.19616, 65.34042, 66.46867, 67.92143, 69.12704, 68.19686, 68.46086,
    69.39777, 66.62844, 60.88995, 59.20912, 61.23245, 52.28214, 53.80286,
    53.74465, 52.50601,
  60.28483, 60.79655, 60.86451, 60.41412, 59.48546, 61.89267, 64.118,
    65.97715, 65.10042, 66.23067, 66.80046, 66.88903, 66.94833, 67.11443,
    66.91278, 66.21336, 66.13585, 67.59987, 69.29012, 70.15026, 70.46187,
    67.39865, 59.72234, 54.81157, 51.51444, 51.93468, 52.15659, 51.28819,
    51.45511, 51.6585,
  60.43167, 59.7477, 61.80385, 62.05518, 62.34986, 62.78855, 63.35177,
    63.73716, 64.40346, 65.03574, 65.74403, 66.27708, 67.04186, 67.59509,
    67.37952, 67.19959, 66.82793, 66.7057, 66.96721, 64.98152, 58.78421,
    58.69827, 55.68736, 52.50274, 53.40459, 52.85607, 52.44907, 51.76181,
    51.05413, 50.99158,
  58.12218, 59.95539, 60.68025, 61.9039, 62.46792, 62.96691, 63.45044,
    63.70608, 63.80685, 64.27351, 65.12924, 66.10012, 67.19541, 68.19736,
    68.30965, 67.96841, 67.91833, 66.80928, 60.27378, 58.04, 55.87237,
    55.43183, 53.70433, 52.73157, 52.68576, 52.5248, 51.99455, 51.44427,
    51.11018, 51.02567,
  62.10343, 60.87752, 61.63078, 62.50019, 63.09291, 63.29545, 63.72457,
    64.04469, 64.04497, 64.02708, 64.34193, 65.38876, 66.97315, 68.07491,
    68.76141, 69.26452, 69.67746, 69.72983, 66.70039, 62.25542, 56.82339,
    55.62385, 54.13565, 53.23922, 53.16718, 52.86884, 51.91491, 51.11379,
    50.82016, 50.9112,
  69.15114, 66.67711, 63.88845, 63.64958, 64.82617, 64.85478, 64.91302,
    65.11121, 65.18657, 64.83544, 64.9006, 65.2384, 65.85366, 66.83238,
    67.76797, 68.87713, 70.06832, 71.34769, 72.20593, 70.49416, 62.49234,
    57.05746, 54.79399, 54.34528, 53.64795, 53.30997, 52.29487, 51.07804,
    50.83135, 50.87201,
  78.3387, 73.85439, 69.11986, 63.72529, 66.31149, 65.85266, 66.10584,
    66.32986, 66.13042, 66.45731, 66.48825, 66.38424, 64.20617, 62.65696,
    61.60332, 63.02422, 67.22375, 70.75694, 72.60252, 73.88713, 70.40581,
    62.36401, 56.91288, 56.35115, 54.874, 54.09801, 52.97069, 51.46796,
    50.82401, 50.92748,
  77.63103, 74.07899, 69.52918, 65.42463, 67.62762, 67.81173, 68.20561,
    68.29355, 68.30057, 68.15111, 68.10532, 67.94238, 68.16293, 66.12507,
    63.18184, 61.81173, 61.94363, 63.88364, 65.5896, 66.39248, 66.64717,
    64.31467, 59.94963, 58.10033, 56.3458, 54.80035, 53.4058, 51.65027,
    50.78599, 50.90586,
  77.93908, 74.40358, 69.85882, 66.49416, 68.80057, 69.08112, 70.20862,
    70.49995, 70.6598, 70.46714, 69.90739, 68.87611, 69.74163, 69.26066,
    67.50539, 66.34904, 65.5151, 65.58475, 65.2199, 63.66682, 62.86775,
    62.73808, 61.80448, 59.71904, 58.10314, 55.94911, 53.90586, 51.8768,
    50.71503, 50.89773,
  77.32982, 74.52661, 69.85417, 67.06654, 69.49413, 70.01595, 71.02052,
    71.90305, 72.70446, 73.25002, 73.22416, 72.62959, 72.28896, 71.91828,
    70.82877, 69.62415, 68.41653, 67.69177, 67.26782, 65.50479, 63.39407,
    62.09133, 62.14444, 60.78584, 59.51846, 56.99052, 54.82105, 52.75382,
    51.04971, 50.83618,
  77.2384, 74.20697, 69.43081, 67.09913, 69.11592, 70.03925, 71.16116,
    72.44146, 74.07852, 75.3045, 75.7868, 76.19579, 76.26644, 76.30092,
    75.97887, 75.63686, 74.53009, 72.98421, 71.1794, 69.17439, 66.6261,
    63.98765, 63.06114, 61.50137, 61.28536, 58.82349, 55.79264, 53.70211,
    52.12416, 51.14923,
  76.68034, 73.4053, 68.70238, 66.35963, 67.90881, 68.82432, 70.50871,
    72.47985, 74.92782, 76.33469, 77.21613, 78.50153, 80.232, 81.21343,
    80.56936, 80.69714, 80.0923, 79.30623, 76.98759, 74.43801, 71.98853,
    68.5747, 65.49098, 63.92424, 63.56792, 61.94612, 58.80171, 54.91034,
    53.37304, 52.06689,
  77.30747, 73.17493, 68.21656, 63.19071, 64.42828, 64.9306, 67.5058,
    71.37186, 73.95394, 74.81747, 76.04413, 77.72498, 79.9576, 80.99141,
    80.63317, 80.82665, 80.44564, 79.13476, 76.9985, 75.65141, 73.44118,
    70.47201, 66.74818, 64.7774, 64.44881, 62.70619, 60.65837, 56.66125,
    53.84698, 52.68282,
  79.2798, 75.41666, 69.54033, 63.29851, 63.10734, 62.63374, 65.0369,
    68.47836, 71.14514, 71.13994, 73.09093, 76.53177, 79.88796, 80.53996,
    78.8507, 78.24924, 77.40156, 75.95547, 74.83521, 74.10291, 72.73846,
    70.38176, 67.29546, 65.31874, 65.34287, 63.81585, 61.81954, 58.40176,
    54.09133, 52.38851,
  80.626, 76.54327, 69.31945, 64.04585, 64.12569, 62.53769, 63.16782,
    64.86458, 65.7458, 66.00343, 67.78772, 71.00525, 74.80119, 75.83846,
    74.3003, 73.37245, 72.27872, 71.47932, 70.84959, 70.94778, 70.35835,
    68.28321, 66.06847, 64.23127, 64.52882, 63.75864, 62.95927, 60.63829,
    55.85848, 52.36194,
  72.14832, 70.94618, 66.38332, 63.80636, 65.1747, 64.45242, 62.88206,
    62.17485, 61.73294, 61.57141, 61.94554, 63.28304, 66.0904, 67.86977,
    67.12292, 66.30263, 65.20521, 64.03297, 64.2728, 65.31727, 65.29671,
    64.23576, 62.00852, 60.57155, 60.56036, 60.06021, 59.51738, 58.68752,
    56.83322, 53.27559,
  57.24886, 58.28507, 59.52409, 60.47913, 61.80437, 63.42484, 61.88538,
    58.4606, 57.33513, 57.65066, 57.09555, 56.85376, 56.82614, 57.49899,
    57.58849, 57.19461, 56.36709, 55.66042, 55.27322, 55.47634, 55.89199,
    56.93726, 57.58948, 57.02179, 56.93684, 56.79087, 56.01954, 54.44,
    53.40618, 52.71768,
  54.39466, 54.61872, 55.13516, 55.22933, 55.85483, 57.615, 58.38862,
    55.85434, 54.35155, 54.84505, 55.09082, 55.11637, 54.85605, 54.42777,
    54.48372, 54.20516, 53.27178, 52.27911, 52.15551, 52.11629, 51.91489,
    52.47881, 53.52727, 54.11043, 53.89745, 53.92987, 53.77386, 52.82629,
    51.79015, 51.165,
  64.69964, 65.34915, 65.87251, 66.52907, 66.86901, 67.01334, 66.72069,
    66.174, 65.60674, 65.28082, 65.22339, 65.27959, 65.26111, 66.23555,
    67.69717, 69.12958, 70.40603, 71.21411, 71.16296, 70.21865, 68.15379,
    65.02451, 62.36884, 60.5835, 58.22952, 54.20705, 51.45513, 53.17315,
    50.73254, 49.07947,
  66.5838, 67.13836, 67.27733, 67.97546, 68.63648, 69.33525, 69.92738,
    69.9575, 69.4934, 68.77647, 67.9589, 67.26978, 66.71352, 66.14303,
    66.01098, 67.03905, 68.88437, 71.56009, 72.18478, 71.8223, 71.34663,
    70.85822, 70.47445, 70.36061, 70.00565, 61.93107, 52.38931, 51.16969,
    50.48578, 49.2824,
  66.89675, 67.60061, 68.32864, 68.74855, 68.6433, 69.05436, 69.93243,
    71.03036, 71.88617, 72.31316, 72.06213, 71.35661, 70.38302, 69.32932,
    68.19691, 66.45959, 65.60845, 66.32649, 68.76947, 71.75069, 71.82219,
    71.77211, 71.60023, 71.29048, 70.53217, 69.34708, 68.47177, 54.65151,
    49.86618, 49.29291,
  67.00744, 67.68948, 68.41363, 69.12914, 69.66465, 70.35394, 70.94289,
    71.20454, 72.3717, 72.70283, 73.14434, 73.95027, 74.36489, 74.15078,
    73.83887, 72.73273, 70.37511, 67.89023, 67.53658, 69.95122, 71.59982,
    71.23642, 67.69934, 70.52949, 69.98649, 70.04451, 69.50714, 68.94746,
    59.06129, 50.75631,
  67.10873, 67.80046, 68.57045, 69.26139, 69.73593, 70.43392, 71.27251,
    71.95133, 72.3446, 72.56716, 73.02375, 74.07152, 74.90982, 74.72375,
    74.47904, 74.37183, 73.81479, 72.97417, 72.24888, 71.44791, 69.65894,
    64.40982, 61.00961, 63.03357, 64.74515, 67.70872, 69.61124, 70.49692,
    70.5583, 60.04441,
  67.22803, 67.88007, 68.68764, 69.41261, 70.00954, 70.79566, 71.90718,
    72.80566, 73.10463, 73.20454, 73.55767, 74.51659, 75.3578, 75.01154,
    74.88832, 74.50746, 73.57642, 73.30915, 72.95211, 72.06805, 71.10892,
    61.02731, 64.93037, 64.19916, 63.67648, 62.75267, 62.86763, 69.54102,
    69.74895, 54.43098,
  67.85819, 68.20896, 68.88209, 69.47768, 70.03479, 70.97131, 72.23456,
    73.30395, 73.9381, 74.0414, 74.28873, 74.24561, 65.93134, 66.63013,
    65.86087, 65.65788, 67.65915, 67.32761, 65.11397, 65.40194, 63.75699,
    63.00681, 65.30555, 67.65931, 67.99358, 67.04613, 67.34264, 69.70843,
    65.44197, 48.19096,
  69.79939, 69.36839, 69.75056, 70.0988, 70.5487, 71.41602, 72.24358,
    67.34963, 62.11288, 64.81465, 65.04078, 64.95989, 65.42976, 66.08451,
    66.46665, 66.49186, 66.09692, 65.38344, 64.30148, 63.29469, 62.74892,
    62.98029, 64.55698, 67.22485, 69.44577, 70.2428, 70.2229, 69.52863,
    61.05339, 48.35334,
  74.1431, 72.7858, 71.96688, 71.72481, 71.74646, 71.93102, 71.41295,
    67.41715, 65.48239, 63.41032, 63.05624, 63.28644, 63.936, 65.76437,
    67.36482, 67.21265, 67.99437, 69.19798, 69.70853, 68.61905, 67.03811,
    66.17181, 65.70551, 65.21228, 67.06726, 70.44654, 70.58133, 68.58042,
    48.37903, 48.93158,
  79.57867, 78.76298, 77.00746, 75.45396, 74.40951, 73.13513, 71.96526,
    72.57929, 72.86259, 69.5387, 65.05379, 63.32291, 62.36344, 61.60691,
    61.49756, 62.57498, 63.8722, 65.31462, 67.10675, 68.61575, 70.33456,
    69.80991, 68.54007, 67.06718, 67.43148, 69.51182, 68.28584, 53.63004,
    48.34456, 48.4022,
  82.52438, 83.08206, 83.88405, 81.80447, 79.67812, 76.39388, 74.50185,
    73.59417, 73.48275, 74.21192, 73.20204, 66.08318, 63.42687, 60.92972,
    59.09743, 58.83676, 58.28345, 58.42351, 59.66946, 61.92632, 65.67924,
    67.35352, 67.78725, 69.70244, 70.34976, 69.89243, 55.74009, 48.91842,
    49.2866, 48.5192,
  80.83102, 81.05315, 85.00952, 86.81776, 85.76556, 81.74534, 77.62132,
    74.40144, 73.35365, 73.84219, 73.58364, 72.97045, 72.80515, 71.64774,
    66.35493, 62.53902, 62.08554, 60.33307, 58.85564, 58.72762, 61.38101,
    63.01976, 62.1687, 65.02553, 69.64704, 69.17328, 48.9539, 53.47688,
    50.1111, 49.05924,
  72.21375, 74.38148, 76.93983, 80.23738, 82.98505, 83.12077, 77.29653,
    73.06799, 75.62987, 74.57883, 74.40507, 73.91994, 74.13105, 74.08697,
    73.2484, 66.5213, 68.7366, 69.40082, 66.8854, 62.37849, 62.92809,
    63.85073, 62.02186, 57.09817, 55.9739, 57.04284, 49.58035, 51.18857,
    50.90466, 49.72755,
  69.83319, 70.35416, 67.64458, 66.32833, 67.31794, 72.41969, 74.27988,
    75.38758, 74.02837, 74.57207, 74.79275, 74.28762, 74.16893, 74.23246,
    73.40453, 72.27411, 71.24184, 71.92075, 71.86423, 70.9157, 65.32893,
    61.30173, 54.29589, 51.14146, 48.8795, 49.08062, 49.18514, 48.70773,
    48.88972, 48.98901,
  70.03508, 66.05019, 67.92113, 67.42601, 67.60986, 68.30733, 70.00806,
    70.47726, 70.8232, 70.38089, 69.94997, 68.29178, 69.95673, 71.0959,
    73.1255, 73.16323, 71.63374, 66.5974, 64.48813, 61.20341, 55.08045,
    55.0732, 52.53001, 49.56381, 50.39135, 50.02779, 49.53712, 48.97884,
    48.40946, 48.4102,
  62.16266, 63.79153, 64.5928, 65.55441, 66.09084, 67.71431, 69.66212,
    71.02644, 70.91997, 70.17691, 70.18722, 70.20576, 70.53747, 71.54649,
    68.52693, 66.73779, 66.43403, 61.22019, 56.88898, 55.07492, 53.25668,
    52.18316, 50.23436, 49.57108, 49.87949, 49.96413, 49.32939, 48.84277,
    48.51883, 48.46228,
  63.79626, 62.76936, 62.98219, 63.33013, 63.45457, 63.67825, 64.72645,
    66.89635, 68.31802, 68.7266, 69.13212, 72.03658, 76.31761, 76.48753,
    72.51889, 70.70571, 68.0796, 64.97231, 60.64336, 57.23408, 53.65073,
    52.63657, 50.80048, 49.84728, 50.09635, 50.0964, 49.21007, 48.5582,
    48.36829, 48.47673,
  70.77406, 67.2628, 64.59444, 63.93507, 63.92191, 63.61706, 63.77021,
    64.32321, 65.33073, 64.94827, 66.12415, 67.85899, 70.1173, 72.44737,
    71.74929, 73.09752, 73.92165, 72.5713, 69.67444, 64.54617, 57.94821,
    53.89891, 51.71749, 50.93088, 50.43248, 50.16068, 49.3849, 48.50583,
    48.42734, 48.46655,
  84.65607, 78.35917, 69.53352, 64.19708, 65.40003, 64.57333, 64.63226,
    64.65025, 64.06207, 64.07228, 64.04676, 63.01536, 61.16317, 60.70612,
    60.79469, 62.93635, 67.30383, 71.78124, 72.63081, 71.29765, 65.53008,
    58.24506, 53.84369, 52.80573, 51.48935, 50.74591, 49.81806, 48.7605,
    48.45082, 48.53413,
  84.5293, 79.23335, 71.33302, 66.50962, 67.48787, 67.06127, 67.02589,
    66.74076, 66.68211, 66.87563, 66.6003, 65.32705, 64.29755, 61.1813,
    58.63309, 57.72736, 58.73716, 61.40265, 63.26065, 63.67805, 63.10966,
    60.11742, 56.35929, 54.46149, 52.75912, 51.4504, 50.19807, 48.90353,
    48.43863, 48.50742,
  85.37074, 81.11997, 72.77864, 68.81866, 69.98597, 69.80947, 70.07446,
    69.91959, 69.70473, 69.14088, 67.68295, 66.37354, 66.48248, 65.35762,
    63.31201, 61.80991, 60.93935, 60.8346, 60.58931, 59.09932, 58.47853,
    58.76448, 58.02338, 55.87321, 54.31526, 52.43433, 50.58251, 49.04686,
    48.38287, 48.50999,
  84.48962, 81.44534, 73.6404, 70.14407, 72.24915, 72.43535, 73.19866,
    73.6181, 74.15845, 73.97781, 72.32827, 70.52087, 69.48535, 68.27899,
    66.81535, 65.31674, 63.68349, 62.73757, 61.71893, 59.70255, 57.42482,
    56.83955, 58.60241, 56.57003, 55.72611, 53.39098, 51.31831, 49.59735,
    48.56815, 48.45264,
  83.06739, 81.0946, 73.73984, 70.14111, 72.78593, 73.74122, 74.86924,
    75.90186, 77.81949, 78.61504, 77.99647, 77.78899, 77.14558, 75.91384,
    73.88442, 72.08212, 70.10314, 68.07953, 66.08051, 63.6574, 60.60109,
    58.44332, 58.90633, 57.2626, 57.31239, 55.02716, 52.38935, 50.50221,
    49.29293, 48.65372,
  82.34333, 79.23607, 73.00298, 70.00183, 71.52654, 72.07949, 74.00497,
    76.32826, 80.05177, 81.41415, 81.08794, 82.87694, 84.72531, 85.02142,
    82.9794, 80.88892, 78.28896, 75.3847, 72.51788, 69.72658, 67.0067,
    64.01277, 60.99472, 59.42229, 59.36361, 58.09736, 55.26619, 51.71111,
    50.35594, 49.33644,
  81.29504, 76.60696, 69.4006, 65.63795, 66.46884, 67.00542, 69.66962,
    74.05737, 78.28941, 78.07781, 77.63419, 79.42899, 82.16515, 83.15399,
    81.73878, 80.62169, 78.51074, 75.8193, 74.04301, 71.84968, 69.12295,
    65.95335, 62.29203, 60.21027, 59.85606, 58.67113, 56.83844, 53.33105,
    50.79259, 49.79298,
  80.99413, 75.94276, 69.35762, 64.61452, 64.30316, 64.03745, 66.43427,
    70.71241, 73.82592, 73.2561, 74.19814, 76.22742, 78.81721, 79.52327,
    78.37589, 77.62904, 75.79358, 73.63497, 72.38688, 71.44101, 68.97004,
    66.28586, 63.05832, 60.94891, 60.90385, 59.31649, 57.60545, 54.24026,
    50.83809, 49.49216,
  77.38646, 73.71184, 67.80815, 63.52895, 63.17161, 61.63256, 62.55382,
    64.67125, 66.24857, 66.35313, 67.90039, 70.29808, 73.17387, 74.30365,
    73.214, 72.3562, 71.1454, 69.41295, 68.82398, 68.43517, 66.70505,
    64.15529, 62.39301, 60.59365, 60.99172, 60.0924, 58.73079, 56.22995,
    51.99108, 49.3864,
  70.14652, 68.67307, 64.48633, 61.92207, 62.8047, 61.91453, 60.71042,
    60.04573, 59.93406, 59.92879, 60.21483, 61.79009, 64.19642, 65.4722,
    65.06969, 64.38899, 63.22721, 62.45853, 62.53625, 63.18269, 62.25498,
    60.43526, 58.31445, 57.32623, 57.60325, 57.30746, 56.40668, 55.26735,
    53.23573, 50.14439,
  56.0144, 56.93602, 57.72107, 58.04243, 59.05533, 60.55295, 58.72933,
    55.79561, 54.87672, 55.01973, 54.42179, 54.04519, 54.23404, 54.71475,
    54.55475, 54.35441, 53.93433, 53.38131, 53.34004, 53.49569, 53.50768,
    54.08697, 54.29834, 53.76842, 53.77436, 53.73515, 53.04482, 51.52021,
    50.67888, 49.96315,
  52.16513, 52.54864, 53.03582, 53.0106, 53.5888, 55.18882, 55.51714,
    53.13267, 51.94951, 52.41946, 52.44515, 52.30349, 52.10534, 51.85093,
    51.60675, 51.38365, 50.57138, 49.80626, 49.80113, 49.81587, 49.65256,
    50.16822, 51.02631, 51.40932, 51.31147, 51.3374, 51.05464, 50.02131,
    49.21571, 48.66356,
  61.20538, 61.31049, 60.89805, 60.51975, 59.9451, 59.52278, 59.16271,
    58.92625, 58.88023, 59.23241, 60.14257, 60.82104, 60.54838, 60.81866,
    60.84822, 60.05927, 58.70816, 57.04987, 54.86373, 52.5194, 50.02454,
    47.39641, 46.19904, 46.30802, 45.80494, 42.6215, 40.42956, 41.9989,
    38.40762, 36.57259,
  65.16186, 65.52637, 65.01088, 64.88018, 64.23553, 63.56884, 62.96605,
    62.22085, 61.39148, 60.76354, 60.70853, 61.24899, 61.97233, 62.2126,
    62.63869, 63.48227, 63.51421, 62.3044, 60.90456, 59.47513, 58.22161,
    57.2161, 56.71126, 56.87793, 56.90901, 51.87466, 38.9575, 40.61623,
    38.39489, 36.93207,
  66.40212, 67.05774, 66.93468, 66.83637, 66.57814, 66.52338, 66.50113,
    66.35601, 65.69776, 64.49488, 63.21964, 62.04076, 60.9045, 60.33843,
    59.87585, 59.16262, 59.8952, 61.86926, 61.31498, 60.2314, 59.49348,
    58.94154, 58.45016, 58.21374, 57.65572, 56.18715, 51.2967, 41.58627,
    37.67036, 37.04621,
  68.07859, 69.19667, 69.44037, 69.74287, 69.53724, 69.47633, 69.57979,
    69.73987, 69.29153, 68.5109, 68.0774, 68.20775, 67.76437, 64.91933,
    63.43013, 61.83447, 59.52338, 58.97477, 61.42878, 60.67878, 59.81249,
    58.67567, 58.0826, 58.26543, 57.68367, 56.79974, 56.08518, 55.30657,
    43.70827, 37.82981,
  68.36467, 70.14753, 70.89036, 71.44414, 71.00188, 70.81039, 70.81306,
    70.18442, 69.20847, 68.07891, 67.69431, 68.42892, 68.71379, 67.8199,
    66.87942, 66.12875, 64.59157, 62.61164, 61.43767, 60.66257, 59.22256,
    53.13071, 52.99844, 57.08562, 57.50098, 57.10907, 56.91337, 57.38904,
    57.04866, 45.99417,
  66.63545, 69.23501, 70.92228, 71.75646, 71.12822, 71.21851, 71.94193,
    71.62276, 70.68219, 69.70249, 69.15716, 69.3524, 69.548, 68.76993,
    68.36694, 67.53836, 65.38013, 63.4165, 61.09967, 59.89117, 58.41356,
    49.32593, 53.04724, 54.53717, 57.13659, 57.26197, 57.47324, 58.08363,
    57.11836, 40.23277,
  65.96576, 67.45942, 69.10405, 70.9546, 71.21542, 71.54075, 72.59566,
    72.76126, 72.06739, 71.04071, 70.10974, 68.83632, 61.73754, 62.20871,
    61.76828, 60.94315, 61.21407, 59.85738, 57.30238, 56.7156, 53.96602,
    52.3318, 53.91444, 56.08205, 57.01767, 56.92629, 57.37904, 57.40276,
    55.01572, 35.69214,
  69.96866, 69.29955, 69.91295, 70.97974, 71.15531, 71.51968, 71.99928,
    68.70827, 64.59456, 66.2635, 65.0758, 63.04319, 61.6839, 61.03476,
    60.32297, 59.74732, 58.96216, 57.33738, 55.14908, 53.78336, 53.34767,
    53.93538, 55.84064, 57.27502, 57.10955, 57.19641, 57.51818, 56.84399,
    46.80056, 35.88331,
  72.63591, 72.25333, 71.57881, 71.27599, 70.84171, 70.51495, 63.24005,
    61.60317, 62.50206, 62.58552, 63.21351, 63.44399, 63.62222, 65.58221,
    66.45456, 64.12473, 63.75616, 63.72816, 62.02829, 58.59463, 55.98987,
    55.75812, 57.20394, 57.03479, 57.08675, 57.66099, 57.30639, 55.04399,
    36.13961, 36.48596,
  75.64413, 75.15432, 73.83144, 72.99713, 72.24559, 70.64314, 62.86234,
    65.29343, 62.06438, 60.09722, 58.53189, 58.93603, 58.84248, 58.62048,
    58.4823, 59.87912, 60.87605, 61.29797, 61.46577, 61.48968, 60.15498,
    58.28996, 56.48174, 56.08843, 56.91849, 57.60038, 56.56136, 41.29768,
    35.90043, 35.82954,
  79.77385, 79.03094, 79.45398, 77.16742, 76.22907, 72.88765, 70.44231,
    68.83195, 67.9905, 67.1106, 58.7127, 53.41662, 52.87464, 51.74664,
    50.79313, 50.77502, 50.95767, 51.4812, 52.75446, 55.22593, 59.60693,
    58.64931, 56.69275, 56.30043, 56.7951, 56.39684, 43.32252, 36.26636,
    36.84204, 35.91697,
  84.1439, 83.2813, 84.80635, 84.96864, 81.87634, 77.69116, 73.56804,
    69.78075, 67.58627, 67.06447, 65.67806, 64.24667, 61.59739, 59.65277,
    56.89452, 52.8325, 52.04575, 50.54527, 49.5287, 50.01667, 53.57233,
    55.61526, 55.28214, 56.68221, 56.81683, 54.49947, 36.69307, 40.79119,
    37.71289, 36.52163,
  76.74905, 78.93229, 80.65464, 82.14792, 82.59164, 80.57105, 73.55214,
    69.04742, 69.93648, 67.88274, 66.62555, 65.50405, 64.9276, 64.74593,
    64.1553, 58.0074, 59.15055, 58.2044, 55.33625, 52.10526, 53.2836,
    54.1115, 51.5573, 46.85812, 46.16866, 44.32242, 37.49472, 39.13143,
    38.80049, 37.2873,
  71.49866, 71.93743, 70.89436, 69.79542, 70.3831, 70.97273, 71.67112,
    71.16849, 68.35352, 68.02412, 67.02975, 65.05073, 64.52396, 64.41018,
    63.29588, 62.48434, 62.12513, 61.37542, 60.74987, 59.17082, 56.48885,
    52.92661, 46.00902, 39.66166, 36.55091, 36.96426, 36.71888, 36.33012,
    36.6691, 36.62449,
  72.04216, 68.54164, 69.03455, 67.31497, 66.21019, 66.06328, 67.52612,
    67.16313, 64.3844, 63.3124, 62.30334, 61.02935, 63.33055, 63.24705,
    63.8744, 63.9099, 62.04971, 60.77752, 58.93204, 55.27084, 48.10944,
    44.57597, 39.76921, 37.78314, 38.28201, 37.72075, 37.08426, 36.5143,
    36.08719, 35.9798,
  64.18171, 67.29707, 68.47387, 69.18195, 69.21167, 70.37148, 71.70374,
    71.15079, 67.9051, 64.2866, 62.75676, 61.42142, 60.83499, 62.1754,
    59.33314, 57.50708, 57.57558, 52.61736, 48.33287, 44.82104, 41.36312,
    40.16734, 38.10184, 37.44696, 37.8222, 37.7288, 36.8908, 36.44614,
    36.15862, 36.02242,
  60.85345, 61.03744, 61.99775, 63.35366, 64.4472, 65.45194, 67.14956,
    69.54617, 70.14974, 68.58231, 66.43175, 67.8743, 68.91339, 68.04021,
    63.21273, 60.49513, 57.6472, 54.92278, 50.81152, 46.70243, 41.98967,
    40.6506, 38.49326, 37.61935, 37.83314, 37.77259, 36.73038, 36.01628,
    35.95534, 35.9673,
  64.81982, 62.57666, 60.62769, 60.47127, 60.99637, 61.60569, 62.83902,
    64.75345, 66.34004, 66.7713, 68.54703, 69.95033, 69.99895, 68.96783,
    67.71286, 67.50606, 66.87181, 64.44031, 60.08643, 53.2381, 45.41301,
    41.6008, 39.40642, 38.54305, 38.02944, 37.61081, 36.82567, 35.94204,
    35.86802, 35.87645,
  79.3627, 72.51761, 63.91065, 58.81701, 59.62002, 58.95705, 59.30555,
    59.75234, 59.71072, 60.37555, 61.42407, 60.86652, 59.14635, 59.11745,
    58.7909, 60.55002, 65.22279, 68.97397, 66.83254, 62.02395, 53.34795,
    45.59327, 41.32636, 40.13403, 38.91119, 38.11398, 37.21148, 36.1746,
    35.82213, 35.90535,
  81.22422, 75.1339, 66.44745, 61.21285, 61.43753, 60.61095, 60.43148,
    60.26239, 60.37919, 60.91021, 60.63923, 58.89089, 58.18856, 55.37985,
    52.64806, 51.7531, 53.18458, 56.33923, 57.21082, 55.45295, 52.62898,
    48.10951, 43.88034, 41.80114, 40.14899, 38.67304, 37.56346, 36.34511,
    35.82036, 35.88656,
  84.52582, 78.94302, 69.90474, 65.02389, 64.99854, 63.92885, 63.51335,
    63.09863, 62.80943, 62.21452, 60.43249, 59.08212, 59.67611, 58.60247,
    56.52097, 54.95496, 54.15987, 53.98646, 53.24617, 50.69238, 48.80314,
    47.72499, 45.67956, 43.59515, 41.40683, 39.34399, 37.78716, 36.43027,
    35.85828, 35.91775,
  85.24226, 82.14536, 73.49206, 69.58729, 70.18376, 69.07839, 68.68929,
    68.05321, 67.79554, 66.47108, 63.70592, 61.72296, 60.9081, 59.77404,
    58.04969, 56.55406, 55.10611, 54.14278, 53.26675, 51.73496, 49.81907,
    47.27397, 45.72813, 44.68397, 43.02135, 40.22338, 38.31331, 37.04771,
    36.05345, 35.86143,
  84.81735, 83.32907, 75.17072, 71.92, 73.67713, 73.72427, 73.54654,
    73.12424, 73.78015, 73.03702, 70.6639, 69.87083, 68.85105, 67.02909,
    64.41518, 62.2544, 59.76651, 56.98323, 54.82597, 52.67601, 50.50425,
    47.89196, 45.70361, 45.072, 44.9627, 42.49306, 39.68573, 38.05687,
    36.82393, 36.03448,
  83.95618, 81.35495, 74.99744, 72.19882, 73.02296, 72.7789, 73.85425,
    75.40508, 78.78713, 78.74261, 77.14639, 78.02307, 78.75905, 78.44278,
    75.65147, 72.78097, 69.25606, 65.18362, 61.23708, 57.46952, 54.04584,
    51.08474, 48.17332, 46.79456, 46.94241, 46.21957, 43.24405, 39.62956,
    38.0892, 36.71345,
  82.39252, 78.01676, 70.82705, 67.52308, 67.50883, 67.31126, 69.92107,
    74.57416, 79.17655, 77.70369, 75.74918, 76.60316, 77.91964, 78.13828,
    76.35647, 74.40855, 71.14964, 67.74727, 65.31721, 61.88335, 57.39894,
    53.50877, 49.66455, 47.3164, 47.33777, 46.85521, 45.34134, 41.61298,
    38.99767, 37.46189,
  80.44568, 76.50729, 70.57124, 66.28362, 65.07497, 64.35228, 67.4144,
    72.46823, 75.61884, 73.9817, 74.21378, 75.14391, 76.42879, 76.48151,
    74.49447, 72.57169, 69.73184, 67.21771, 65.50516, 63.0896, 59.50777,
    55.41898, 51.51511, 49.12805, 48.83544, 47.76436, 46.25834, 42.78662,
    38.74669, 37.05361,
  76.40928, 73.01096, 67.43051, 63.45835, 62.61755, 60.8251, 62.22462,
    65.12897, 66.93137, 66.65027, 68.078, 69.82416, 71.59161, 71.78949,
    69.69209, 67.5814, 65.44532, 63.54001, 62.24217, 60.53023, 57.46021,
    54.89661, 52.15363, 50.43929, 50.436, 49.76501, 48.61137, 45.57737,
    40.24761, 36.72289,
  68.27818, 65.94996, 62.4747, 59.66729, 59.96195, 58.76756, 57.70321,
    57.16215, 56.33847, 56.56887, 57.06187, 58.35944, 60.17997, 60.66544,
    59.72253, 58.48165, 56.84246, 55.73384, 55.61618, 55.07204, 52.87238,
    49.85352, 47.31358, 46.21235, 46.59936, 46.51791, 45.93328, 45.05372,
    42.59425, 37.93109,
  51.47956, 52.19141, 52.38702, 52.36332, 53.12494, 54.56669, 52.11716,
    48.13894, 46.85274, 46.98759, 46.46671, 46.00786, 45.95003, 46.1279,
    45.9068, 45.70824, 44.7951, 44.05627, 43.67093, 43.27755, 42.76822,
    42.86558, 42.57933, 41.9489, 42.11663, 42.17676, 41.46911, 39.98735,
    39.13902, 37.86514,
  43.57615, 44.04123, 44.25595, 43.85828, 44.35849, 46.22407, 46.58902,
    43.0661, 41.29723, 41.9254, 42.21286, 42.28025, 41.95161, 41.46391,
    41.09921, 40.7414, 39.47501, 38.22682, 38.02369, 38.00796, 37.74223,
    38.18758, 38.9901, 39.31981, 39.12015, 39.38591, 39.22185, 37.92747,
    36.86957, 36.09555,
  49.35227, 49.21763, 49.12418, 49.15928, 49.0134, 49.12305, 49.40566,
    49.73927, 50.18676, 50.90231, 52.01453, 51.83155, 49.57277, 49.34169,
    49.19201, 48.47458, 48.09073, 48.02258, 47.90237, 48.10008, 47.54561,
    45.80387, 45.91824, 47.57756, 48.31462, 46.43244, 47.24768, 48.54966,
    39.02156, 35.57641,
  53.82572, 53.48746, 52.41314, 52.4664, 51.7067, 51.39165, 51.80661,
    52.33583, 53.15039, 54.23846, 55.7192, 57.67617, 59.05589, 58.24426,
    57.87109, 58.57647, 58.20728, 58.99624, 59.89275, 60.46749, 59.97249,
    58.94489, 58.48775, 60.67797, 62.21518, 53.14299, 43.4445, 46.10884,
    39.15402, 36.47006,
  56.16673, 56.06316, 55.66162, 55.04666, 54.31963, 53.89816, 53.67175,
    53.59916, 53.70846, 53.94967, 54.52147, 55.70452, 57.2154, 59.1484,
    60.55925, 60.04251, 61.20063, 61.98458, 62.71369, 63.43081, 64.14371,
    64.68073, 64.80774, 64.77552, 64.21416, 62.47897, 53.36319, 45.25273,
    38.30016, 36.89701,
  59.89817, 60.21814, 60.59809, 60.2035, 59.76466, 59.5012, 59.29571,
    59.12804, 59.11119, 59.02173, 59.02094, 59.53766, 59.26273, 58.31554,
    60.33574, 61.59983, 60.02265, 59.47973, 62.31718, 63.38167, 64.40341,
    64.77582, 65.17625, 65.76098, 65.13231, 63.82035, 62.2114, 53.18671,
    42.34568, 36.6985,
  61.90156, 61.22709, 60.9192, 60.40596, 59.78197, 59.45793, 59.40179,
    59.22112, 59.25769, 59.2592, 59.42223, 60.2305, 60.93998, 61.24918,
    61.80732, 62.59484, 62.52528, 61.75024, 62.04359, 63.07586, 63.53133,
    58.73565, 59.97453, 64.81486, 65.19402, 64.3167, 62.88639, 62.96082,
    62.67432, 44.61574,
  62.02472, 61.7504, 61.61543, 61.17982, 60.26982, 60.01334, 60.46088,
    60.1381, 59.6003, 59.44263, 59.77636, 60.7501, 61.85308, 62.23102,
    63.32267, 64.49645, 64.44978, 63.55715, 62.63864, 63.03869, 61.68054,
    53.73439, 58.54724, 61.99305, 64.47936, 64.1314, 63.4832, 64.03268,
    62.9288, 40.01253,
  62.06749, 61.91843, 61.87856, 61.56899, 60.94299, 60.98559, 61.72553,
    61.67588, 61.1458, 60.71509, 60.5446, 60.30257, 60.07867, 60.80673,
    61.76619, 62.83067, 63.38307, 62.80795, 59.91667, 60.43928, 58.25826,
    57.51754, 60.28082, 63.84325, 64.17531, 61.90929, 63.57847, 63.38486,
    56.67888, 34.47043,
  62.22402, 62.07907, 62.19603, 62.1035, 61.80201, 62.14937, 62.62328,
    61.55813, 60.82838, 61.02563, 61.02364, 61.13737, 61.4517, 62.07137,
    62.72819, 63.4858, 64.12836, 63.97507, 60.52297, 59.74467, 60.31368,
    62.65592, 65.13991, 65.33387, 64.43159, 64.05096, 64.39707, 63.43074,
    50.05246, 35.2357,
  63.33081, 62.9407, 62.47225, 61.96343, 61.2962, 61.26227, 61.0537,
    61.64497, 62.17447, 62.60268, 62.98342, 63.16201, 63.60841, 65.23453,
    66.25125, 65.28551, 65.77766, 66.493, 66.42046, 65.45329, 63.99803,
    65.37249, 66.23571, 65.90073, 64.90384, 65.41846, 64.42403, 59.49442,
    37.40001, 35.79909,
  64.69181, 65.05848, 63.96377, 63.70773, 62.69637, 61.20656, 59.92874,
    60.75342, 61.02733, 61.8386, 62.65281, 63.27547, 63.19, 63.19801,
    63.30273, 64.70913, 65.51685, 65.98382, 66.30794, 66.81551, 67.07066,
    65.68378, 64.01528, 60.23755, 63.69379, 64.36898, 62.87719, 43.87894,
    35.1991, 33.98723,
  64.72013, 64.48322, 65.73376, 64.31168, 64.80772, 62.8821, 61.94761,
    61.69915, 62.20196, 62.88028, 61.62315, 52.36576, 49.92737, 50.23283,
    50.47446, 52.1565, 53.8346, 55.15273, 57.04083, 61.761, 66.58627,
    65.71265, 59.29908, 59.49267, 62.49952, 59.4629, 43.73941, 35.68614,
    35.93699, 34.19324,
  70.31045, 68.5065, 70.17069, 70.78322, 68.39709, 65.95584, 63.69247,
    61.33295, 59.88559, 60.19901, 60.10057, 59.69528, 60.45253, 60.86756,
    53.37136, 52.92632, 52.06189, 51.82205, 52.06562, 54.9037, 61.9738,
    63.58311, 58.22772, 63.14991, 62.84983, 54.09082, 36.43011, 40.33009,
    37.15308, 35.21207,
  69.15173, 70.61571, 72.24586, 73.35284, 73.04418, 70.65364, 63.85097,
    60.5274, 62.31529, 61.05202, 61.3938, 61.3336, 62.50266, 63.13725,
    61.93716, 58.94592, 58.64658, 58.14437, 56.2109, 57.0632, 59.641,
    58.51487, 54.499, 50.49613, 49.30209, 45.28163, 37.33486, 39.02784,
    38.74077, 36.31671,
  61.09513, 61.21919, 61.6292, 60.98844, 60.94188, 61.41763, 62.66483,
    63.09354, 61.38938, 62.06726, 62.78022, 62.62623, 63.96403, 64.57775,
    63.41824, 62.16164, 61.92536, 62.87096, 63.64286, 63.57301, 59.31601,
    54.88041, 48.16201, 41.39025, 37.86372, 37.38494, 36.09985, 35.45874,
    35.90642, 35.48892,
  63.99705, 63.72537, 62.49182, 61.38868, 60.8377, 61.34101, 63.0234,
    63.19667, 61.53913, 61.74827, 61.74491, 61.38652, 61.94785, 62.89441,
    62.7968, 61.95675, 62.04399, 62.99155, 64.24522, 61.85193, 50.20154,
    47.02729, 41.15413, 39.16147, 39.2902, 37.98206, 36.6278, 35.71758,
    34.93673, 34.52731,
  64.5404, 64.82378, 64.52538, 63.65875, 62.92503, 63.24771, 63.83373,
    63.37588, 62.22897, 61.35269, 61.33967, 60.87704, 59.46634, 61.63293,
    60.81045, 60.13321, 60.9364, 57.2887, 55.62179, 50.806, 43.34797,
    43.03655, 39.36632, 38.36026, 38.71034, 38.08594, 36.25882, 35.79577,
    35.10443, 34.58931,
  60.42159, 60.33831, 61.76886, 62.71312, 62.6782, 62.45057, 62.80832,
    63.61423, 63.48846, 62.79688, 61.90181, 62.72514, 63.99838, 63.29877,
    62.10638, 60.72305, 57.89687, 56.52762, 55.93353, 51.83411, 42.99547,
    43.1762, 40.00922, 38.47804, 38.35206, 38.01752, 35.93016, 34.71062,
    34.58212, 34.43724,
  58.24152, 57.59033, 56.43734, 57.98486, 59.7793, 61.83094, 62.17138,
    62.89466, 63.45535, 63.32569, 64.26635, 65.32175, 65.58327, 65.90256,
    65.3028, 65.0137, 65.27396, 66.05435, 64.68085, 56.73714, 44.96654,
    42.56705, 40.28654, 39.23859, 37.6807, 36.77871, 35.96379, 34.39399,
    34.28437, 34.17966,
  69.47363, 63.26431, 55.44712, 51.67029, 53.53596, 54.06932, 55.702,
    57.62141, 58.60015, 61.04583, 62.86527, 63.01997, 60.52605, 63.29297,
    64.33474, 65.62112, 68.36032, 70.83439, 70.75658, 68.78124, 55.66197,
    46.9456, 42.3677, 40.47106, 38.1647, 36.8338, 35.92386, 34.7162,
    34.25198, 34.20869,
  68.80988, 63.02912, 55.39904, 50.70372, 51.52452, 51.69703, 52.57253,
    53.74582, 55.76055, 59.23229, 59.56702, 54.69366, 54.93042, 53.86647,
    52.67654, 52.82952, 56.47109, 62.32233, 65.24943, 63.9661, 59.28608,
    52.82066, 46.54037, 42.82682, 40.11959, 37.58933, 36.23891, 34.90586,
    34.23509, 34.22163,
  70.32516, 65.15543, 57.07587, 52.31067, 52.10294, 51.62998, 51.95269,
    52.72218, 54.25174, 55.61357, 53.01919, 50.1656, 53.19646, 53.19876,
    51.8967, 51.19935, 51.92017, 53.34108, 54.89579, 54.25973, 54.23658,
    54.94981, 52.04778, 47.13349, 42.38755, 38.7052, 36.45966, 35.04713,
    34.27593, 34.22596,
  74.48525, 70.28551, 62.89411, 59.07246, 58.77291, 56.88797, 56.52856,
    56.13252, 57.52268, 56.89231, 52.21977, 50.07483, 51.54363, 51.66567,
    51.03176, 50.92466, 50.3255, 50.46802, 51.50314, 52.20593, 52.87172,
    52.58614, 52.47959, 51.6039, 47.15929, 40.51992, 37.32909, 35.91877,
    34.51926, 34.18984,
  77.26745, 75.97185, 69.20086, 66.04284, 67.6104, 67.09326, 65.65565,
    63.63011, 64.01075, 62.01822, 57.52362, 58.03654, 58.28935, 57.84503,
    56.22925, 55.88748, 54.52044, 51.6841, 50.71705, 50.60179, 50.37834,
    49.48473, 48.86128, 50.10089, 50.8553, 45.3859, 39.86198, 37.77752,
    35.86731, 34.41449,
  77.4707, 76.02298, 71.90314, 69.70485, 69.71432, 68.83566, 69.34568,
    69.83539, 72.49664, 70.87312, 66.40726, 68.95275, 70.69479, 70.8294,
    68.88774, 66.88755, 64.17712, 60.44055, 56.73446, 54.43072, 52.60334,
    50.90134, 49.43699, 49.48846, 51.07162, 51.30627, 46.47056, 40.3334,
    37.98481, 35.4984,
  76.78519, 73.55678, 68.62453, 64.89558, 64.59707, 63.82001, 65.74924,
    70.61681, 73.93877, 71.88721, 66.81587, 69.44255, 71.23835, 71.93003,
    70.99409, 70.25182, 68.0708, 65.85881, 63.50149, 60.48902, 57.29345,
    54.2892, 51.19194, 49.39772, 50.07159, 51.24701, 50.53681, 44.38738,
    39.98878, 37.29188,
  75.62953, 72.77291, 68.6431, 65.88764, 63.13487, 61.68993, 65.89089,
    70.75674, 72.73605, 68.82063, 68.29099, 69.83536, 71.68663, 71.51419,
    69.87655, 68.86305, 67.97646, 67.23194, 66.63514, 65.16747, 63.10986,
    60.25662, 56.15469, 53.41165, 53.2243, 52.19384, 51.4437, 46.11946,
    38.38942, 36.07246,
  72.37697, 69.93667, 66.76859, 64.36144, 62.27402, 59.46421, 61.97369,
    64.96778, 65.03186, 63.43339, 65.39662, 67.3511, 68.90546, 69.23917,
    67.82565, 65.82615, 64.70084, 64.76222, 64.89073, 64.34817, 63.26586,
    62.8633, 61.70733, 59.76249, 59.68393, 59.1214, 58.79379, 54.03141,
    42.1161, 35.18823,
  67.67653, 66.22816, 64.07309, 63.08645, 63.80718, 63.7312, 61.80266,
    59.21876, 56.22838, 57.11124, 58.06352, 59.8672, 61.71906, 62.45354,
    62.34779, 60.91014, 59.06466, 58.68268, 59.50885, 60.2094, 58.04349,
    54.35349, 51.76181, 51.51727, 52.87337, 53.72719, 54.01818, 55.21499,
    50.37896, 38.656,
  55.89629, 56.77118, 57.50648, 58.56322, 62.05723, 63.64629, 61.24183,
    52.95758, 50.7225, 51.74504, 51.02726, 50.72478, 51.31105, 52.05293,
    52.38304, 51.95183, 50.48859, 49.39335, 48.11768, 46.21146, 45.40002,
    44.77564, 43.62949, 42.8996, 43.98336, 44.93694, 44.79935, 42.60499,
    41.94778, 39.10992,
  47.595, 48.17742, 48.19102, 47.89056, 50.15478, 55.34723, 56.67879,
    48.56487, 45.1052, 47.77273, 49.30298, 50.0494, 49.84574, 49.06909,
    47.75486, 46.38507, 42.81124, 39.64604, 39.3275, 38.8619, 37.66362,
    38.07201, 38.64293, 39.08833, 39.40894, 40.40936, 40.46915, 38.34685,
    35.96584, 34.25488,
  41.42599, 41.59044, 41.67392, 41.81453, 41.76808, 42.03923, 42.4941,
    43.07581, 43.79227, 44.86383, 47.24211, 47.11768, 43.12993, 43.42859,
    43.93266, 43.43158, 43.59467, 44.62526, 45.78261, 47.71095, 48.40336,
    46.68866, 47.40644, 50.26826, 52.35223, 51.98208, 57.3342, 59.07917,
    43.43269, 39.47011,
  45.12518, 45.54137, 44.61061, 45.51555, 44.83526, 44.46128, 45.12216,
    45.84069, 46.5974, 47.58091, 49.23742, 51.4525, 52.46703, 49.8298,
    48.33135, 49.19254, 48.1896, 49.34077, 51.32714, 52.92657, 52.32609,
    51.4, 51.98771, 56.02967, 58.59313, 54.76118, 52.35941, 56.99231,
    44.91162, 40.8913,
  43.87166, 44.49495, 45.40179, 46.19197, 46.85429, 47.33736, 47.47802,
    47.93073, 48.51932, 49.24927, 50.3121, 51.82576, 53.30938, 55.42305,
    56.60235, 54.49384, 54.80992, 56.45836, 57.51075, 58.63834, 58.89088,
    59.05033, 59.15227, 59.64195, 59.55129, 58.39925, 58.17269, 54.92552,
    44.64114, 42.28153,
  47.0509, 47.6656, 49.42929, 51.23122, 52.75169, 54.25385, 54.1729,
    53.42558, 53.8852, 54.71555, 54.94524, 55.80622, 55.50681, 54.32444,
    57.95601, 60.43316, 57.58053, 54.71658, 57.81376, 59.04784, 59.46848,
    59.62315, 60.12701, 61.15848, 61.27027, 60.30886, 58.62033, 55.15595,
    46.21878, 40.56952,
  49.74664, 49.16627, 51.41651, 53.12278, 54.46968, 54.66259, 54.61621,
    54.47295, 55.88251, 57.05238, 57.18744, 59.69678, 60.85973, 60.6586,
    60.72184, 61.19574, 60.43213, 57.14923, 58.38829, 58.98579, 59.01358,
    57.06992, 58.84243, 60.59454, 61.71495, 60.74669, 58.26366, 58.01514,
    58.04485, 46.43169,
  51.72453, 54.27071, 58.19529, 61.77582, 61.65911, 61.73296, 62.49266,
    62.36134, 61.59242, 61.18517, 61.14902, 61.6325, 62.13092, 61.75266,
    62.16016, 62.87247, 62.27282, 60.44768, 58.65135, 58.8131, 58.50942,
    53.99947, 58.26052, 60.10808, 61.08878, 60.39251, 58.6929, 59.0727,
    58.59504, 44.53322,
  52.66392, 55.42029, 59.12437, 61.90826, 61.58615, 61.62135, 62.00903,
    61.79118, 61.14369, 60.94509, 60.92556, 60.90975, 59.97833, 61.36295,
    61.72614, 61.94738, 62.04094, 60.65873, 58.66734, 59.1686, 58.31178,
    57.52114, 59.64387, 60.91861, 60.92991, 59.3236, 58.96647, 58.85416,
    58.06974, 39.83987,
  52.89343, 55.58268, 59.5279, 62.53927, 62.37936, 62.43058, 62.89309,
    61.59554, 55.74873, 57.16733, 57.50084, 57.90805, 58.92885, 62.11634,
    62.54758, 62.85072, 63.29182, 62.73771, 61.08471, 60.58319, 60.13496,
    60.32327, 61.34158, 61.89033, 60.74337, 59.8199, 60.16723, 59.62015,
    56.15204, 40.29771,
  63.16729, 63.81568, 64.24516, 64.06406, 62.99193, 62.9119, 63.12087,
    63.56701, 64.27498, 64.59654, 64.67511, 64.94345, 65.66244, 68.36747,
    69.62441, 66.59442, 66.67966, 67.16241, 66.44846, 64.16193, 62.55194,
    63.43383, 64.90565, 64.09097, 61.88786, 62.43019, 61.2014, 59.32222,
    44.90411, 39.92478,
  68.90769, 70.36226, 69.65319, 70.13207, 68.17393, 65.92478, 64.37838,
    65.11162, 65.5247, 67.14445, 68.21264, 68.9061, 68.22004, 66.61001,
    64.98767, 66.22559, 66.52739, 66.26648, 65.92443, 66.61738, 66.98593,
    64.85331, 63.19045, 61.00642, 60.62414, 60.73644, 59.56192, 49.28651,
    40.01274, 37.06313,
  67.31925, 67.24696, 68.77211, 68.21234, 68.56866, 66.96225, 65.63658,
    65.37184, 65.90678, 65.90497, 63.66212, 56.94978, 55.62888, 55.97509,
    57.12106, 59.14861, 60.62597, 61.09179, 61.90818, 62.76266, 64.29578,
    63.4971, 59.25907, 57.02238, 57.85415, 57.76315, 46.97278, 40.03556,
    39.45206, 37.23883,
  72.35606, 70.50279, 73.728, 74.24458, 71.58698, 68.56406, 66.01895,
    63.29272, 60.91236, 58.50115, 54.9693, 53.07895, 56.0325, 58.11748,
    57.63523, 56.8327, 55.94592, 56.69038, 58.30038, 60.65605, 63.16703,
    62.66013, 58.67308, 58.95379, 58.45757, 52.50343, 40.79034, 42.79116,
    40.9681, 38.40697,
  76.43578, 78.39114, 80.17211, 79.97009, 78.32458, 74.19782, 65.94549,
    62.15801, 62.85984, 60.5655, 60.5636, 59.83085, 60.63777, 61.38282,
    60.98489, 60.09222, 60.26892, 60.42599, 61.23533, 62.95484, 62.46443,
    61.13853, 57.55893, 55.64381, 54.71114, 48.85937, 42.02177, 42.95709,
    43.01785, 39.81422,
  67.49776, 68.28441, 68.73335, 67.45454, 66.81714, 67.72771, 69.23876,
    68.91848, 65.22237, 64.59634, 64.16702, 61.94981, 62.88892, 63.4332,
    61.72499, 60.39688, 60.1332, 60.20616, 60.71092, 60.97471, 59.95684,
    55.96082, 52.61961, 48.52077, 44.49902, 43.39735, 40.69144, 39.55975,
    40.08197, 39.04749,
  64.46078, 65.35931, 65.79263, 65.7171, 65.22493, 65.82397, 68.63016,
    68.50629, 65.26824, 64.09499, 62.75582, 61.93146, 62.59996, 62.77267,
    61.90687, 61.18807, 60.57958, 61.07141, 62.15432, 61.47701, 50.86639,
    51.56561, 47.76869, 46.16972, 45.48288, 43.26983, 41.2508, 39.59293,
    38.53854, 37.78084,
  65.2102, 65.8082, 66.2616, 65.87169, 65.28413, 65.99508, 67.04625,
    65.98104, 64.24359, 62.97012, 62.90872, 61.54358, 60.74412, 62.09039,
    61.43068, 61.04367, 61.49271, 61.53169, 62.20753, 60.88264, 48.5084,
    48.79807, 44.81387, 44.17757, 44.53399, 43.32046, 40.54056, 39.63785,
    38.75825, 37.87066,
  59.09032, 56.7216, 58.50262, 61.27715, 64.16848, 63.83746, 64.3026,
    65.60648, 65.02711, 63.96932, 62.28289, 62.98584, 65.25476, 63.6206,
    61.55294, 61.25283, 61.09657, 61.18451, 62.09346, 61.15224, 47.50781,
    49.04766, 45.57072, 43.8331, 43.00356, 42.44476, 40.05621, 38.23137,
    38.02262, 37.65999,
  55.66819, 56.61766, 56.82994, 59.57859, 62.46964, 64.18227, 63.71331,
    63.77039, 64.20998, 63.24633, 64.35989, 66.19956, 65.59818, 64.21677,
    64.37417, 63.04073, 62.00545, 62.59465, 63.75916, 61.26816, 48.7267,
    47.10001, 45.28327, 44.66028, 42.22523, 40.81767, 39.9496, 37.56628,
    37.49252, 37.28764,
  61.01173, 58.03603, 53.58285, 51.90614, 54.18465, 55.78202, 57.47494,
    58.53349, 58.75224, 62.21318, 63.68406, 63.16032, 60.13812, 61.62981,
    62.1764, 62.97158, 65.21985, 67.53751, 68.21413, 65.57508, 59.14109,
    50.18163, 46.07208, 44.34732, 41.42715, 39.92579, 39.22437, 37.87798,
    37.4277, 37.25544,
  60.17357, 57.91643, 53.16343, 50.67884, 52.09287, 53.06109, 53.9868,
    55.35442, 58.55452, 64.03591, 64.24622, 60.30065, 59.37946, 58.36761,
    57.41264, 57.89957, 61.5954, 63.44592, 64.23248, 63.82967, 61.86959,
    57.1463, 49.94096, 46.60101, 43.87503, 40.75086, 39.4079, 37.96426,
    37.38953, 37.24783,
  58.36158, 56.68933, 51.47809, 48.69652, 49.18576, 49.94131, 50.84443,
    52.31344, 56.02709, 61.32952, 58.68798, 53.57806, 57.97619, 57.91663,
    56.23883, 54.50032, 55.22103, 56.24747, 57.66961, 58.77443, 59.57472,
    60.97152, 57.5665, 52.08337, 46.41906, 41.91063, 39.32086, 38.19504,
    37.53936, 37.3134,
  57.46965, 53.42925, 50.59527, 49.39297, 49.70478, 48.55138, 49.67417,
    50.90618, 55.81982, 58.01682, 51.45928, 47.4628, 50.80145, 52.03615,
    52.12236, 52.86727, 53.19618, 53.81015, 55.3991, 56.07313, 56.68188,
    57.99594, 59.74854, 58.63811, 51.54728, 43.35002, 39.67563, 39.002,
    37.82206, 37.30429,
  58.18904, 57.30894, 53.52837, 52.77019, 55.95394, 57.15544, 56.10498,
    54.07674, 56.18084, 54.84386, 48.07852, 48.94497, 51.16922, 52.87922,
    52.75323, 54.53298, 55.07048, 52.44804, 51.7977, 51.84408, 51.32336,
    51.31425, 51.73467, 54.47078, 56.56095, 49.72116, 43.08714, 41.19297,
    39.55364, 37.54045,
  65.71255, 64.95695, 60.99482, 60.29538, 61.04728, 60.38108, 62.25191,
    63.28196, 66.4295, 60.7595, 52.65483, 55.06229, 57.41517, 59.77611,
    59.57457, 59.79417, 60.02874, 57.98321, 54.51964, 52.84593, 51.2442,
    50.09827, 49.97084, 50.40561, 53.51096, 56.77793, 51.94299, 43.62519,
    41.44495, 38.59571,
  67.95004, 65.15403, 58.64166, 56.6132, 58.67192, 59.17079, 59.78579,
    63.09221, 69.06651, 64.82356, 55.94003, 57.98063, 59.09372, 60.39804,
    60.89421, 62.71796, 63.07034, 62.85346, 60.15255, 56.47956, 54.21007,
    52.86716, 51.3476, 49.78373, 51.09174, 55.94653, 57.16322, 50.19685,
    45.5037, 41.37886,
  72.81381, 71.52899, 67.93774, 61.33536, 59.41428, 59.34448, 64.29693,
    68.18275, 67.11148, 61.30157, 60.35681, 61.77943, 62.123, 61.78368,
    61.29244, 63.25086, 65.67821, 67.0105, 66.19841, 64.12749, 62.0156,
    60.68754, 57.64485, 54.50678, 54.38608, 55.04827, 57.32841, 52.41891,
    43.59763, 40.20716,
  72.53059, 71.10417, 65.81665, 61.518, 60.3292, 58.15633, 63.21192,
    65.71621, 61.89741, 60.10097, 62.1319, 61.95952, 61.87708, 62.34488,
    63.42192, 65.02192, 67.1885, 67.47129, 67.03399, 66.36999, 65.67329,
    65.63617, 65.17674, 64.37936, 63.77999, 62.93831, 62.5139, 61.01945,
    46.96677, 38.10466,
  66.34261, 67.18987, 66.4528, 66.81219, 68.18722, 67.40118, 65.94393,
    62.01966, 55.92479, 58.01633, 59.12438, 59.38991, 59.69167, 60.78131,
    63.1913, 63.88837, 63.70108, 65.41278, 65.66755, 65.54049, 64.37327,
    62.7818, 60.70419, 60.34653, 61.57013, 61.98473, 61.86794, 62.03778,
    60.39082, 42.59167,
  60.01213, 61.07287, 63.61219, 65.39561, 66.867, 68.38103, 67.69167,
    59.42154, 55.46634, 56.70033, 56.20542, 57.80759, 59.39093, 59.72066,
    61.02339, 61.41185, 59.85797, 58.74036, 55.65661, 51.5281, 50.90453,
    49.32106, 46.17392, 45.35255, 47.20486, 49.51336, 50.2261, 48.81723,
    48.70133, 43.90477,
  57.35953, 58.42434, 59.47138, 60.08349, 64.18791, 66.73441, 67.20242,
    62.13834, 56.21538, 60.11134, 63.02813, 63.60535, 63.16406, 61.74019,
    59.86456, 57.68775, 52.04884, 46.90864, 46.017, 44.53038, 42.3952,
    42.30229, 42.23742, 42.23143, 43.02284, 44.83084, 45.43551, 42.99005,
    39.74871, 37.27728,
  38.60357, 39.08539, 39.52832, 39.99334, 40.364, 40.81763, 41.34529,
    41.92015, 42.54474, 43.29611, 44.88314, 45.00932, 43.04637, 43.51556,
    43.77676, 43.33695, 43.42921, 43.92051, 44.52144, 45.81307, 46.42664,
    45.68906, 46.23182, 47.46467, 48.13157, 47.57819, 50.61509, 50.6391,
    40.66449, 37.44546,
  44.51176, 45.31709, 45.38976, 46.56148, 46.87605, 47.34793, 48.21135,
    49.02008, 49.89952, 50.78838, 51.78735, 53.02576, 53.65845, 52.27477,
    51.58248, 51.79442, 50.76764, 51.03014, 51.78832, 52.35998, 51.94016,
    51.18421, 51.25054, 53.49766, 57.245, 55.51591, 51.59657, 52.26971,
    41.76656, 38.5499,
  47.33109, 48.42472, 49.45122, 50.67139, 51.8194, 52.96507, 54.0534,
    55.27581, 56.49801, 57.52104, 58.39666, 59.4954, 60.48755, 61.78183,
    62.60624, 61.07483, 60.89602, 61.3087, 61.16939, 61.62903, 62.95022,
    64.0944, 63.79869, 64.01193, 65.56998, 63.08083, 57.10472, 50.98169,
    42.04581, 39.66599,
  52.93966, 54.7602, 56.64819, 58.60426, 60.04557, 60.36023, 60.57867,
    60.67203, 60.82632, 60.80403, 60.84606, 61.44477, 61.93405, 62.16541,
    63.67421, 65.71664, 67.13023, 65.23201, 65.68343, 66.44939, 68.87957,
    67.7364, 63.78002, 67.9925, 69.36838, 63.6653, 59.45877, 49.59151,
    42.08416, 38.17858,
  57.68885, 58.82158, 60.35112, 60.51971, 60.48817, 60.70422, 61.1068,
    61.25949, 61.43268, 61.34378, 61.40211, 62.0764, 62.66101, 63.1466,
    64.10706, 65.979, 67.59084, 64.81303, 64.344, 69.01319, 70.53054,
    62.81718, 62.21058, 64.52044, 67.27277, 65.1508, 58.55724, 58.32594,
    53.86664, 41.50161,
  60.91331, 61.06026, 61.38441, 61.46006, 61.04292, 61.05341, 61.67802,
    61.76946, 61.51765, 61.47868, 61.75875, 62.65876, 63.54486, 63.7775,
    64.61636, 66.67814, 69.35575, 70.38392, 69.0935, 68.42256, 64.46227,
    60.17014, 60.9737, 62.29949, 64.61317, 62.60361, 60.11849, 68.65066,
    61.7927, 40.05641,
  61.5665, 61.59036, 61.81373, 61.74537, 61.25773, 61.28521, 61.80484,
    61.85328, 61.44206, 61.40887, 61.6189, 61.88251, 62.13963, 62.66489,
    63.37729, 65.36424, 68.39275, 68.49181, 63.17006, 62.63722, 60.50623,
    58.96228, 59.5921, 62.00604, 61.50994, 57.63613, 60.43444, 66.78191,
    56.25843, 37.42802,
  61.78703, 61.71795, 61.83094, 61.83671, 61.37999, 61.30682, 61.69921,
    61.35938, 60.88867, 60.98865, 61.22297, 61.47186, 61.72937, 62.24277,
    63.35768, 65.72135, 68.34628, 66.36982, 61.6959, 60.72239, 59.60659,
    59.55415, 61.54764, 62.78707, 59.59994, 58.1908, 64.66039, 62.69177,
    47.4438, 37.84322,
  63.87582, 63.86755, 63.99841, 63.83813, 63.34919, 63.48366, 63.65355,
    64.07903, 64.65915, 64.86691, 65.08195, 65.38963, 65.78718, 67.40482,
    68.99815, 69.27177, 71.61769, 73.9547, 74.54161, 72.88505, 69.40133,
    72.17418, 73.5124, 72.66527, 65.18458, 64.71268, 63.8004, 54.92664,
    41.50417, 37.62394,
  70.12441, 70.36538, 70.34502, 70.70219, 69.64387, 67.90717, 67.3202,
    68.02114, 68.35747, 68.95208, 69.36942, 70.14706, 70.0968, 69.46934,
    69.72726, 72.21584, 74.15768, 74.80759, 74.18009, 72.57681, 71.61349,
    68.61423, 65.99203, 61.03915, 64.81438, 71.1346, 60.7711, 42.40314,
    37.69135, 36.02704,
  71.28465, 71.5382, 73.05812, 72.90588, 73.85618, 72.56059, 71.24417,
    70.70376, 70.34444, 70.56609, 70.05049, 65.25335, 64.68211, 64.98093,
    66.42079, 68.86433, 71.28841, 69.99424, 65.87878, 63.07016, 63.85686,
    59.49308, 51.96045, 48.22211, 49.49785, 48.6698, 42.09576, 37.42923,
    36.9331, 35.97639,
  72.58437, 69.0445, 71.57546, 72.97394, 72.39953, 70.89252, 69.89432,
    67.29005, 64.52029, 64.179, 63.43533, 62.41039, 62.57385, 63.17147,
    64.02281, 66.10131, 63.1653, 60.46258, 57.87941, 56.78509, 57.75451,
    53.69535, 46.60994, 52.02675, 54.58232, 42.49044, 37.41117, 37.99733,
    37.41875, 36.43344,
  79.17288, 79.09073, 80.23271, 80.86206, 79.70406, 75.98277, 68.2342,
    64.65305, 65.62959, 63.38184, 64.01576, 63.41677, 63.56728, 63.9579,
    64.27466, 65.78915, 66.07719, 62.70632, 59.79491, 60.63384, 58.68332,
    51.20395, 47.43787, 48.34023, 48.75172, 41.00021, 38.18874, 38.33883,
    38.29534, 37.0127,
  72.77045, 72.75835, 72.59295, 70.78741, 69.45222, 68.53283, 68.31204,
    68.92252, 66.68932, 66.51551, 67.35873, 65.74816, 66.88107, 67.48309,
    66.37137, 66.6478, 68.69469, 70.84531, 71.63888, 67.46005, 57.66744,
    51.46722, 50.97348, 43.47591, 40.00759, 39.20311, 37.83118, 37.20196,
    37.35973, 36.76694,
  65.41176, 65.06369, 64.83192, 64.45949, 64.51817, 65.85696, 69.5538,
    70.62669, 68.17675, 68.10156, 67.46204, 66.69544, 66.57568, 66.28112,
    66.05831, 66.2822, 68.33041, 70.5402, 71.62898, 66.8838, 53.45685,
    49.32608, 42.85187, 40.50858, 39.26252, 38.72253, 37.75768, 37.02145,
    36.63762, 36.27438,
  66.63836, 66.92923, 67.29843, 67.20287, 67.1595, 68.02912, 68.994,
    68.81841, 68.15789, 67.48518, 66.97298, 65.29826, 64.44753, 65.03726,
    64.71394, 65.95776, 68.51324, 64.30096, 60.71717, 55.97313, 45.11158,
    43.75411, 41.07746, 40.12303, 39.38993, 38.54808, 37.66883, 37.12234,
    36.68493, 36.24895,
  66.28667, 66.02834, 66.0854, 66.19741, 66.71947, 66.64612, 67.116,
    67.74719, 67.26175, 66.65433, 65.44812, 65.4852, 66.31531, 64.8472,
    64.41073, 65.9605, 65.89922, 60.01297, 60.10701, 57.13243, 43.71545,
    43.67907, 41.5361, 40.24598, 39.13757, 38.58505, 37.4575, 36.58207,
    36.41096, 36.19022,
  64.29682, 64.58627, 64.5593, 64.85318, 64.9632, 65.33028, 65.50188,
    65.88721, 66.27644, 65.49774, 65.67072, 66.03803, 65.29224, 64.83262,
    65.46165, 66.43817, 60.69854, 55.8947, 58.0017, 54.01255, 43.96967,
    42.8746, 41.04377, 39.85886, 38.15849, 37.67819, 37.2368, 36.27973,
    36.17202, 36.03323,
  66.12141, 65.0606, 63.88301, 63.14088, 63.5998, 63.61985, 64.02506,
    64.60111, 64.5328, 64.51666, 65.07829, 64.64133, 63.60851, 64.52544,
    65.95038, 68.80357, 72.56593, 73.38363, 73.50612, 66.6234, 52.68553,
    44.5606, 40.77519, 39.60402, 37.65543, 37.14292, 36.86763, 36.33661,
    36.13182, 36.01834,
  65.78426, 64.54679, 63.31831, 62.48176, 63.0549, 63.46859, 63.94707,
    64.32122, 64.63363, 65.32587, 65.35365, 64.10173, 64.07759, 64.58405,
    65.94386, 68.4628, 69.33173, 68.79989, 67.16988, 64.10159, 56.50448,
    48.20752, 42.15585, 40.23656, 38.53352, 37.42559, 36.87562, 36.4174,
    36.13514, 36.02187,
  65.1804, 64.09032, 62.66421, 61.83572, 62.29651, 62.74525, 63.12663,
    63.39977, 63.71117, 64.10408, 63.49748, 62.46797, 62.7147, 63.15995,
    62.60317, 59.50324, 57.70495, 56.70013, 56.7739, 55.51717, 53.42069,
    51.31131, 46.52355, 42.44577, 39.63839, 37.99051, 36.88082, 36.45557,
    36.16027, 36.03033,
  65.45921, 63.58159, 62.30074, 61.38828, 61.59871, 61.63044, 61.85434,
    61.91239, 62.35098, 62.39355, 59.96643, 57.12344, 57.54404, 56.51456,
    54.88216, 53.37226, 51.81123, 50.76656, 50.26314, 49.43838, 50.25737,
    51.09511, 49.61515, 48.36545, 43.71984, 39.10604, 37.07939, 36.75758,
    36.23905, 36.04151,
  65.31033, 63.36941, 61.55376, 61.06634, 61.53654, 61.57543, 61.26852,
    59.91342, 60.13744, 58.03603, 53.77911, 53.88974, 54.27617, 54.01917,
    52.80965, 52.35453, 51.26342, 48.67623, 47.37732, 46.76029, 47.50136,
    48.26131, 46.37583, 46.77293, 46.30828, 41.64978, 38.0345, 37.66033,
    36.84429, 36.12685,
  67.10429, 65.73263, 64.54274, 63.77456, 63.69349, 63.40086, 63.54792,
    63.87727, 64.26268, 61.154, 57.25927, 58.89724, 59.4755, 59.17585,
    57.52935, 55.76208, 54.26885, 51.73491, 48.58738, 47.53164, 47.79134,
    47.36333, 45.76301, 44.72967, 44.93179, 44.69671, 41.24266, 38.33441,
    37.45173, 36.44846,
  69.11095, 69.25296, 66.72404, 65.64848, 65.83403, 65.67893, 65.56831,
    66.10358, 67.12057, 65.56133, 61.15, 62.64801, 62.67215, 61.2905,
    59.11082, 57.22617, 54.7245, 52.79612, 49.97828, 47.32933, 47.1447,
    46.6766, 45.10659, 43.76302, 42.65879, 43.58726, 43.63751, 40.77277,
    38.99004, 37.44061,
  71.83035, 72.1953, 70.07025, 68.47762, 67.89145, 67.46348, 67.93246,
    68.67242, 68.43117, 65.86963, 64.05738, 64.5761, 64.19272, 61.25,
    57.89714, 55.91253, 54.10311, 52.59489, 50.4825, 48.10081, 47.95145,
    47.50526, 45.17425, 43.34331, 42.80766, 43.02124, 43.99547, 42.20294,
    38.76288, 37.2218,
  72.32476, 72.38742, 70.29591, 68.9422, 68.6972, 68.22701, 68.46793,
    68.64555, 67.7011, 64.97845, 64.93587, 64.8211, 63.69029, 61.24147,
    58.96187, 56.94384, 55.22722, 54.37182, 53.01667, 51.67057, 52.98793,
    54.68531, 53.49051, 49.99004, 47.57439, 46.78672, 47.35891, 45.80723,
    39.58638, 36.26306,
  72.52719, 72.33619, 70.82316, 70.16273, 70.52124, 70.1149, 69.51051,
    68.86388, 67.82244, 67.8029, 67.71762, 67.69877, 66.85981, 65.10279,
    64.05311, 62.24745, 59.9557, 58.99852, 58.40843, 58.11089, 58.29999,
    56.66521, 53.1223, 50.50179, 48.83295, 48.05867, 47.14312, 48.41539,
    45.51134, 38.09427,
  68.15193, 67.97874, 68.85715, 69.33292, 69.69814, 69.95626, 68.96977,
    67.15131, 66.43324, 66.49478, 66.18436, 65.8122, 65.6827, 66.54678,
    67.83862, 66.00206, 63.43113, 61.13533, 57.44696, 53.53963, 51.93201,
    49.897, 47.53788, 45.85673, 45.38641, 45.10603, 44.1835, 42.48946,
    41.87619, 39.12197,
  66.95077, 66.8102, 67.19984, 67.21543, 67.73479, 68.83523, 68.73746,
    66.83851, 65.74222, 66.04011, 66.12633, 65.91719, 65.60238, 65.87408,
    65.93681, 61.64789, 56.05479, 51.05705, 48.72232, 46.39946, 44.4515,
    43.53684, 42.74012, 42.04213, 41.6178, 41.61402, 41.13911, 39.48404,
    37.59403, 36.22831,
  34.08419, 34.17002, 34.25272, 34.35608, 34.36852, 34.42526, 34.54763,
    34.69285, 34.87423, 35.12888, 36.07743, 36.26342, 34.85266, 35.06684,
    35.2542, 34.8669, 34.87712, 35.1436, 35.45746, 36.31064, 36.87857,
    36.3506, 36.54885, 37.52808, 38.32715, 38.19016, 40.78988, 42.40994,
    36.7067, 34.85278,
  35.71509, 35.95407, 35.69712, 36.11237, 36.03538, 35.98618, 36.23267,
    36.4686, 36.724, 37.04644, 37.49401, 38.17657, 38.59684, 37.66507,
    37.09459, 37.38897, 36.93317, 37.35152, 38.19326, 38.96212, 39.0788,
    39.00409, 39.56787, 41.02573, 45.70899, 47.02631, 41.03535, 43.41306,
    37.39849, 35.51315,
  37.1843, 37.40748, 37.54726, 37.795, 37.96385, 38.18085, 38.41955,
    38.68795, 38.98212, 39.26418, 39.61542, 40.20546, 40.62745, 41.20835,
    41.51659, 40.62083, 40.80524, 41.64666, 42.08327, 42.86584, 44.38734,
    46.20087, 47.14464, 46.80627, 50.72481, 53.11932, 44.17276, 42.56004,
    37.35913, 36.18631,
  40.50776, 41.03582, 41.64912, 42.31639, 42.96364, 43.81333, 44.10358,
    43.94854, 44.17234, 44.68188, 45.02911, 45.53804, 45.51143, 44.90185,
    46.05896, 47.22026, 46.30104, 44.98149, 45.84402, 46.84856, 49.35189,
    50.10146, 47.75571, 52.52405, 55.01374, 47.92472, 47.06757, 41.65292,
    37.35358, 35.26515,
  45.39448, 45.55047, 46.2674, 46.98511, 47.44732, 47.66548, 47.7688,
    47.83247, 48.46669, 49.1094, 49.02534, 49.16404, 49.1785, 49.41508,
    49.48653, 49.62827, 48.68015, 46.93034, 47.05141, 51.90992, 54.09095,
    45.74806, 45.7213, 47.23378, 49.03245, 47.92567, 44.08718, 44.25615,
    43.65836, 37.39143,
  48.83598, 49.71457, 50.84585, 52.2939, 52.37966, 52.0822, 52.66806,
    53.03691, 53.05457, 53.78684, 54.8089, 57.22523, 59.65643, 58.62074,
    57.45523, 65.34827, 74.76511, 59.89338, 49.59653, 50.24594, 47.66729,
    44.13085, 44.92509, 46.15402, 48.47716, 47.18056, 50.0028, 65.82068,
    57.30629, 36.17977,
  53.50191, 55.18866, 56.85099, 58.70629, 59.55854, 60.28437, 61.87539,
    63.6192, 63.32766, 62.37522, 61.67157, 59.48047, 56.36076, 55.42264,
    59.44735, 65.38806, 59.634, 51.14898, 47.27646, 46.79915, 45.29932,
    44.33279, 44.96985, 47.25224, 48.10237, 44.52679, 54.00164, 71.33615,
    54.67878, 34.34661,
  58.83081, 60.75677, 62.40311, 63.8393, 63.40467, 64.52129, 65.42749,
    60.63105, 56.72548, 55.51839, 53.88267, 51.94601, 50.07066, 49.54939,
    49.69242, 49.89589, 49.34586, 48.09678, 45.11514, 44.52345, 43.78839,
    43.61015, 45.13641, 46.97788, 45.98093, 43.91619, 54.74334, 60.47319,
    41.22526, 35.06177,
  62.69152, 63.1675, 63.66309, 62.96529, 61.25659, 60.90669, 57.39646,
    54.73133, 54.50099, 54.03297, 53.27142, 52.33703, 51.81213, 55.03865,
    56.98452, 51.14366, 50.03881, 51.2427, 50.72456, 47.5889, 45.34521,
    47.56348, 51.78469, 51.92255, 47.17282, 47.66256, 50.51242, 47.23341,
    37.49949, 34.99891,
  68.93815, 70.82469, 70.15317, 70.24093, 67.4175, 61.58765, 55.67168,
    56.94858, 57.42722, 59.0754, 61.09896, 64.35, 64.12228, 60.54124,
    56.51596, 56.98462, 57.26617, 56.4662, 54.30356, 52.92551, 53.24884,
    52.45654, 51.60734, 47.86331, 55.6063, 69.76418, 55.23893, 38.38771,
    35.30354, 33.95325,
  73.47791, 73.61662, 74.54168, 74.07507, 74.10592, 73.7608, 73.03918,
    73.37545, 73.89468, 75.48044, 76.71164, 62.72421, 57.8014, 56.53237,
    55.68722, 55.44948, 55.49238, 54.47866, 52.82018, 51.86248, 53.38198,
    51.16728, 45.85653, 42.42129, 44.29418, 45.66011, 39.64264, 34.93643,
    34.49162, 33.85801,
  78.33507, 75.00156, 78.48062, 80.14738, 80.16135, 78.81982, 77.76348,
    74.86276, 71.7457, 70.97679, 67.22739, 59.25772, 60.77677, 60.21592,
    54.82929, 54.00147, 51.64394, 50.25122, 48.62955, 47.87144, 49.03165,
    46.75941, 40.80586, 45.04501, 47.95283, 37.71172, 34.6404, 35.04299,
    34.80312, 34.1494,
  85.1676, 85.72365, 88.47651, 89.66867, 88.7165, 84.50591, 76.44361,
    72.17313, 72.60668, 70.8182, 71.13011, 66.24748, 67.55261, 67.50617,
    57.61543, 52.43939, 50.07044, 48.44159, 46.77519, 47.79521, 47.74134,
    43.45314, 40.12789, 43.49129, 45.62663, 36.68005, 35.15298, 35.30214,
    35.39243, 34.568,
  82.5396, 84.08748, 83.87154, 81.99197, 79.86421, 77.9426, 76.89063,
    76.83979, 74.41412, 73.25573, 74.27892, 73.26853, 74.89105, 76.96693,
    78.90028, 62.02315, 51.28613, 52.12251, 52.18642, 50.93653, 46.04243,
    44.91357, 47.91034, 40.16739, 36.99694, 36.00528, 35.12101, 34.71448,
    34.8582, 34.43098,
  74.4959, 74.11732, 73.53279, 72.55536, 71.80902, 73.59128, 78.91405,
    79.03761, 75.55643, 74.7309, 73.54033, 72.47944, 70.84041, 73.62064,
    73.82514, 57.40081, 55.33041, 52.91499, 53.49975, 54.65751, 50.87245,
    44.20942, 38.60371, 36.62145, 35.83554, 35.81238, 35.12794, 34.57046,
    34.3182, 34.07658,
  70.97167, 71.18769, 71.75194, 71.87119, 71.96133, 72.89439, 73.91946,
    73.61565, 72.69128, 71.75636, 71.4465, 65.86367, 61.39127, 61.42514,
    57.85048, 54.4425, 52.85682, 49.1336, 47.911, 46.42139, 40.13841,
    38.30093, 36.36521, 35.99622, 35.95118, 35.62532, 35.09282, 34.63561,
    34.32084, 34.04948,
  70.34279, 70.62711, 71.08426, 71.3931, 71.78802, 71.42123, 71.55078,
    72.08483, 69.89655, 67.68145, 62.95397, 62.3408, 64.45085, 58.98586,
    54.4122, 51.68116, 48.92547, 45.84525, 46.62364, 45.73249, 37.54486,
    37.82719, 36.85352, 36.11256, 35.71252, 35.67093, 35.00896, 34.33215,
    34.193, 34.03046,
  69.55558, 69.80627, 68.09613, 67.27725, 66.10474, 65.62991, 65.02077,
    64.47926, 64.14539, 61.41037, 61.5065, 62.939, 60.0709, 57.53473,
    56.45888, 51.21888, 45.54598, 42.6027, 44.86196, 43.79364, 37.80996,
    37.66491, 36.88156, 36.22603, 35.2934, 35.09541, 34.80928, 34.13972,
    34.01633, 33.91707,
  67.82909, 66.2545, 63.01271, 60.89981, 60.19403, 59.27035, 58.78109,
    58.55332, 57.45522, 56.43815, 57.51807, 55.74254, 50.44905, 50.2631,
    49.991, 48.61413, 48.80055, 49.59135, 51.91641, 50.92233, 43.96296,
    39.18679, 36.76862, 36.22527, 35.00989, 34.66017, 34.48679, 34.12869,
    33.98064, 33.90032,
  63.75075, 61.78121, 58.85144, 56.31779, 55.59126, 54.92862, 54.36264,
    53.79548, 53.39595, 54.85719, 54.86171, 50.37271, 48.85149, 48.69999,
    48.29448, 47.63436, 48.58298, 49.8684, 50.44381, 50.14855, 46.34646,
    41.21278, 37.17041, 36.41548, 35.4255, 34.77686, 34.48327, 34.18213,
    33.97935, 33.90034,
  59.97571, 58.30067, 55.52165, 53.32952, 52.47146, 51.98328, 51.59026,
    51.36908, 51.85818, 53.45218, 51.96877, 48.72134, 49.51744, 49.25016,
    47.90925, 46.1453, 45.24636, 44.59242, 44.45552, 43.71788, 42.44468,
    41.45803, 39.36829, 37.50841, 36.02164, 35.12228, 34.50214, 34.19925,
    33.9972, 33.90931,
  59.44731, 56.52137, 54.30396, 52.74452, 52.03614, 51.0553, 50.9233,
    50.76484, 52.14706, 52.79671, 49.73449, 47.52482, 47.58302, 46.42115,
    44.67278, 43.1637, 41.75994, 40.80486, 40.38602, 39.64585, 40.84692,
    41.98284, 40.22305, 40.69762, 38.34817, 35.8019, 34.58432, 34.35038,
    34.03091, 33.92031,
  58.38223, 56.65075, 54.22376, 52.78257, 53.0792, 52.92406, 51.9267,
    50.44741, 50.65544, 49.50436, 46.0016, 45.10069, 44.54425, 43.56612,
    42.03945, 41.48775, 41.02692, 39.57443, 38.85754, 38.41087, 39.52374,
    40.41981, 38.2248, 39.29396, 39.54403, 37.07384, 34.99522, 34.86186,
    34.39625, 33.97287,
  58.54757, 57.20646, 56.02159, 55.28811, 54.66762, 53.46613, 52.94638,
    51.92505, 51.65268, 48.37407, 44.60024, 44.692, 44.54121, 44.10989,
    43.05787, 42.3063, 41.89967, 40.78784, 39.12653, 38.45199, 38.54771,
    38.47313, 37.77934, 37.64373, 38.28907, 38.60175, 36.86876, 35.25867,
    34.79508, 34.18126,
  57.96096, 58.1428, 55.2735, 53.84226, 53.64688, 52.70633, 51.32144,
    50.56495, 51.1899, 48.61594, 44.58571, 45.08432, 45.15306, 44.54477,
    43.58598, 42.95931, 42.00627, 41.44082, 40.20495, 38.77872, 38.70952,
    38.78928, 38.25092, 37.45066, 36.86063, 37.86096, 38.19437, 36.62549,
    35.69259, 34.77606,
  58.52921, 59.91285, 58.22905, 55.38568, 53.51489, 52.27192, 52.68773,
    53.01146, 50.84586, 47.84229, 46.10435, 46.33729, 46.33942, 44.87976,
    43.15356, 42.39447, 41.81664, 41.4591, 40.62658, 39.23055, 39.16583,
    39.12433, 37.96564, 37.02192, 36.91704, 37.375, 38.42918, 37.64961,
    35.66069, 34.65367,
  59.38956, 59.90411, 56.62719, 54.51097, 53.43017, 51.9938, 52.56423,
    52.10832, 49.08302, 46.82708, 46.62437, 46.5482, 45.93596, 44.42031,
    43.04738, 42.04354, 41.27227, 41.08024, 40.46003, 39.372, 39.89161,
    41.40411, 41.65594, 40.18991, 39.32258, 39.31344, 40.32072, 39.91839,
    36.12385, 34.04482,
  58.8903, 58.15004, 55.99939, 55.15576, 54.74937, 53.39226, 52.61637,
    50.59304, 47.08261, 46.41487, 46.04143, 45.81183, 45.24179, 44.08389,
    43.57674, 42.7636, 41.74809, 41.79099, 42.16899, 42.43794, 43.19575,
    43.28888, 41.92945, 40.74107, 40.07605, 40.04796, 39.90422, 41.26955,
    39.79903, 35.22881,
  56.56669, 55.29959, 55.52706, 56.00488, 55.58343, 55.53398, 53.14332,
    48.51764, 45.99725, 45.85025, 44.92124, 44.35965, 44.17731, 44.29829,
    44.96289, 45.17747, 44.99247, 45.04827, 43.98064, 42.27901, 41.808,
    41.02513, 39.75971, 38.90089, 38.84065, 38.95732, 38.63935, 37.94344,
    37.90255, 35.96931,
  55.84742, 55.62657, 55.15182, 54.18682, 53.85857, 55.42612, 55.30714,
    50.29758, 47.1496, 48.02373, 48.58728, 48.97263, 48.75535, 48.37587,
    47.91544, 46.88525, 44.77743, 42.40946, 41.26046, 39.94076, 38.85631,
    38.33516, 37.86965, 37.47174, 37.26386, 37.36264, 37.09446, 36.1389,
    35.14012, 34.16996,
  28.64926, 28.69121, 28.72995, 28.77149, 28.76688, 28.77472, 28.8068,
    28.86938, 28.97005, 29.11433, 29.87471, 30.08723, 29.02993, 29.18609,
    29.32039, 28.97436, 28.91432, 29.0092, 29.10868, 29.68305, 30.04891,
    29.5111, 29.51031, 30.15174, 30.68888, 30.59654, 32.96043, 34.65787,
    30.73605, 29.37972,
  29.25637, 29.37374, 29.09992, 29.37762, 29.24362, 29.12875, 29.25238,
    29.37678, 29.50937, 29.7064, 30.07265, 30.60234, 30.96704, 30.31421,
    29.84178, 30.00761, 29.53586, 29.7044, 30.26099, 30.80822, 30.79637,
    30.5202, 30.88308, 31.92916, 36.35747, 38.3068, 33.52542, 36.05095,
    31.38055, 29.88729,
  29.428, 29.45606, 29.45026, 29.51105, 29.52001, 29.56063, 29.64429,
    29.7833, 29.91711, 30.03485, 30.21687, 30.64456, 30.96587, 31.44334,
    31.71314, 30.94135, 30.97996, 31.57485, 31.83291, 32.32824, 33.47047,
    34.98988, 36.13176, 35.9554, 40.64433, 44.22564, 35.72479, 35.28319,
    31.22769, 30.41582,
  30.29191, 30.40132, 30.65842, 30.95262, 31.28841, 31.83554, 32.0017,
    31.8111, 31.90339, 32.21401, 32.36461, 32.69677, 32.69059, 32.30796,
    33.38946, 34.55473, 34.11098, 33.23817, 33.96854, 34.87495, 37.2471,
    38.51266, 36.92439, 41.80317, 44.92623, 38.59499, 38.08136, 34.25078,
    31.18492, 29.73274,
  32.53733, 32.42788, 32.87904, 33.34681, 33.6846, 33.83958, 33.92883,
    33.93183, 34.3869, 34.81393, 34.59828, 34.57301, 34.55952, 34.93052,
    35.57347, 36.24649, 35.81376, 35.20749, 35.75932, 40.64156, 43.15024,
    35.99564, 35.85754, 37.34812, 38.97035, 37.94218, 35.34423, 35.2126,
    35.48995, 31.32604,
  34.715, 35.21184, 36.027, 37.06793, 37.00028, 36.53493, 36.8742, 37.071,
    36.96669, 37.37465, 37.90975, 39.6753, 41.7016, 41.47816, 40.73635,
    48.60255, 58.7038, 46.7952, 38.60099, 39.94257, 38.05849, 34.55667,
    34.95033, 35.67892, 37.6647, 36.92331, 39.64039, 54.11508, 48.44631,
    30.50363,
  37.34837, 38.25298, 39.27871, 40.51048, 41.0186, 41.46393, 42.93625,
    44.94019, 45.41733, 45.43316, 45.70724, 44.61338, 42.50118, 41.72132,
    46.92595, 55.15447, 49.79363, 40.56627, 37.43487, 36.97161, 35.50562,
    34.54875, 34.9224, 36.6627, 37.82236, 35.04835, 44.48854, 62.54828,
    47.84559, 29.00007,
  40.78629, 42.26502, 43.87106, 45.59803, 46.05921, 48.02307, 50.24477,
    47.89832, 45.63225, 45.20237, 44.08011, 42.16966, 40.04347, 39.13652,
    39.69565, 40.528, 39.27376, 37.88679, 35.7518, 35.26324, 34.61153,
    34.28712, 35.41032, 37.02047, 36.65801, 34.63084, 46.7174, 54.49465,
    34.93585, 29.95816,
  46.5867, 47.8751, 49.11557, 49.56863, 49.32304, 50.0622, 48.0389, 45.90392,
    45.38843, 44.55464, 43.14998, 41.4462, 40.03717, 42.0717, 43.57522,
    39.16101, 38.47359, 39.67555, 39.32011, 36.79488, 34.87183, 36.43274,
    39.96331, 40.35327, 36.67416, 37.14747, 41.2896, 40.18932, 32.21605,
    29.88987,
  52.70094, 55.03746, 55.35236, 55.6907, 54.11639, 49.77573, 44.72021,
    44.77597, 44.33765, 44.44292, 45.27034, 47.87135, 47.66264, 45.10168,
    42.06026, 41.94495, 42.24047, 41.885, 40.59965, 40.13034, 40.5415,
    40.90771, 41.29211, 38.72663, 46.32045, 59.20881, 46.95905, 32.8264,
    30.2897, 28.81345,
  74.72932, 77.03868, 69.52872, 60.31926, 58.17114, 55.07214, 51.15265,
    53.1292, 54.62046, 62.72049, 69.99424, 48.31798, 42.47873, 40.98626,
    39.91992, 40.22683, 41.5765, 41.20719, 40.21983, 39.91516, 42.39525,
    41.60679, 37.70807, 34.91678, 38.21191, 41.27681, 35.0561, 29.85086,
    29.30173, 28.66857,
  86.63454, 79.34652, 84.82259, 86.9578, 82.95399, 70.24012, 70.4488,
    64.01896, 53.39996, 55.97833, 54.63587, 42.37816, 43.74981, 43.86448,
    39.59139, 40.57532, 39.39531, 38.82964, 38.02824, 38.02499, 40.35547,
    38.92236, 33.81863, 37.37748, 39.80186, 31.99225, 29.26626, 29.67752,
    29.55437, 28.93835,
  89.8833, 90.93419, 95.69202, 97.54394, 97.71123, 94.88776, 79.33713,
    55.6879, 56.23805, 51.49908, 50.09407, 44.37204, 47.59248, 48.60199,
    41.35886, 40.6172, 39.47599, 38.29047, 37.08945, 38.86742, 39.96845,
    36.12465, 33.07637, 37.29245, 39.34385, 31.06548, 29.62657, 29.84995,
    30.08609, 29.32749,
  91.93094, 97.49784, 97.58027, 95.66197, 92.93612, 89.26443, 85.6493,
    85.82806, 76.22789, 72.29253, 80.48663, 76.09552, 75.81403, 72.8932,
    62.72398, 48.39413, 39.84251, 41.34413, 42.24503, 42.43026, 38.80917,
    37.57858, 40.09432, 34.37213, 31.64158, 30.39433, 29.68271, 29.35124,
    29.65481, 29.24833,
  80.41494, 80.17127, 74.66127, 70.37058, 65.87791, 76.80122, 88.14137,
    89.05351, 86.64388, 85.82987, 82.02312, 64.03909, 51.37446, 56.25107,
    60.69274, 44.42122, 44.10344, 43.29361, 46.08916, 47.79689, 42.68782,
    37.78526, 33.33572, 31.0091, 30.11285, 30.39423, 29.77969, 29.29868,
    29.13016, 28.87953,
  64.11707, 61.955, 61.02964, 60.06448, 60.73998, 65.2515, 70.02282,
    67.38615, 63.95595, 60.01135, 54.99689, 48.35341, 44.86588, 46.85464,
    45.75389, 43.25442, 43.87656, 41.47976, 41.90474, 41.55125, 34.98727,
    32.33505, 30.39546, 30.27953, 30.52365, 30.30033, 29.8036, 29.38008,
    29.10568, 28.83501,
  59.60165, 58.08165, 57.3432, 57.23746, 57.70233, 57.31447, 56.45244,
    55.67467, 53.59586, 50.94864, 46.66992, 46.84575, 50.24634, 46.36111,
    43.11885, 42.31182, 40.86529, 38.38067, 40.18291, 39.73661, 31.41334,
    31.53153, 30.99327, 30.46562, 30.26303, 30.31058, 29.74918, 29.09884,
    28.97085, 28.81724,
  55.73378, 55.50416, 54.39743, 53.90777, 52.9805, 52.34426, 51.75449,
    51.09679, 49.95297, 47.62257, 47.3156, 49.39149, 47.48492, 45.80685,
    46.59563, 43.1734, 38.03847, 35.08846, 38.17416, 37.76914, 31.68297,
    31.81616, 31.38404, 30.82845, 29.84126, 29.82304, 29.57487, 28.89744,
    28.78291, 28.70717,
  55.18027, 54.1548, 51.59929, 49.7441, 48.98471, 48.20494, 47.77031,
    47.6134, 46.56094, 45.42234, 46.76853, 45.28604, 39.60036, 39.45591,
    39.86739, 38.67607, 38.54293, 39.10537, 42.17722, 42.04288, 36.13013,
    33.04993, 31.57021, 30.91109, 29.67979, 29.41888, 29.29081, 28.90811,
    28.74476, 28.68235,
  52.94656, 51.37469, 48.92668, 46.88627, 46.35878, 45.9088, 45.53674,
    45.06402, 44.45119, 45.58598, 45.15713, 39.52362, 36.53218, 36.13457,
    35.91952, 35.39418, 36.7554, 38.80336, 40.86675, 41.8701, 39.00119,
    35.04296, 31.8694, 31.01988, 30.07659, 29.47504, 29.24581, 28.94948,
    28.7547, 28.69752,
  49.98695, 49.00727, 47.17736, 45.27923, 44.59067, 44.1537, 43.58825,
    42.90958, 42.79711, 43.76467, 40.94996, 35.93794, 35.89358, 36.02182,
    35.73013, 34.96065, 34.97376, 35.3167, 36.33782, 36.666, 36.07253,
    35.55333, 33.80849, 31.83472, 30.47954, 29.76338, 29.24796, 28.96756,
    28.77531, 28.69354,
  48.97002, 47.65396, 45.64897, 44.27283, 43.48386, 42.28098, 41.7795,
    41.16219, 42.14568, 42.30992, 38.18126, 35.20538, 35.52737, 35.36029,
    34.86197, 34.33979, 33.65099, 33.2158, 33.16665, 32.7348, 34.2395,
    35.39406, 34.44156, 35.11331, 33.01118, 30.544, 29.36128, 29.11525,
    28.82545, 28.71402,
  47.88232, 46.31702, 43.99974, 42.60216, 42.87667, 42.91852, 42.26009,
    41.20605, 41.9435, 40.69772, 36.43111, 35.03009, 34.74952, 34.45196,
    33.77314, 33.87693, 33.70491, 32.42198, 31.76253, 31.52381, 33.14059,
    33.97392, 32.28165, 33.88963, 34.32869, 31.77021, 29.66645, 29.61794,
    29.17134, 28.75354,
  46.81496, 45.2258, 44.27621, 43.87109, 43.78692, 43.54764, 44.04766,
    44.08603, 44.66005, 41.10951, 36.09053, 35.37434, 35.04634, 35.00576,
    34.61696, 34.45712, 34.51551, 33.56492, 32.02246, 31.67887, 32.18077,
    32.28351, 31.66026, 31.82774, 32.85955, 33.22104, 31.45503, 29.99932,
    29.54979, 28.94515,
  46.22238, 46.71378, 44.2742, 43.38843, 43.92171, 43.9572, 43.44855,
    43.55646, 44.74756, 41.34792, 35.97073, 35.39735, 35.20636, 35.04831,
    34.81092, 34.82706, 34.46808, 34.23635, 33.05516, 31.65738, 31.93502,
    32.34439, 32.13868, 31.35876, 30.73194, 31.98196, 32.3924, 31.04517,
    30.42621, 29.49964,
  47.22362, 48.98581, 47.89815, 45.90598, 44.50773, 43.49769, 44.41252,
    45.51802, 43.5772, 39.70713, 36.59389, 36.04229, 36.0479, 35.15573,
    34.2386, 34.08849, 33.97372, 34.13774, 33.4751, 32.02832, 32.40017,
    32.79479, 31.6908, 30.72319, 30.49693, 31.05871, 32.42151, 31.89342,
    30.37467, 29.42697,
  48.69087, 49.86419, 46.86404, 44.95266, 43.98076, 42.77469, 44.03854,
    44.38521, 41.17987, 38.02082, 36.72114, 36.07691, 35.64631, 34.74884,
    34.11839, 33.76507, 33.53281, 33.74469, 33.21887, 31.92699, 32.63792,
    34.54813, 34.90028, 33.29867, 32.37857, 32.51171, 34.07826, 34.10424,
    30.69859, 28.83498,
  48.20607, 47.88906, 45.77361, 44.99789, 45.03311, 44.13945, 44.3086,
    42.80686, 38.92324, 37.53938, 36.35412, 35.63824, 35.13345, 34.48864,
    34.57518, 34.21202, 33.45287, 33.56792, 33.84037, 33.76849, 35.17896,
    36.16761, 35.03268, 33.67535, 32.94463, 33.17949, 33.44115, 35.42865,
    34.13144, 29.84124,
  45.49987, 44.29378, 44.59882, 45.78308, 46.38852, 47.19199, 45.47091,
    41.26402, 38.42616, 37.50125, 35.49967, 34.02733, 33.36219, 33.67032,
    34.83841, 35.42025, 35.59466, 36.08602, 35.19793, 33.64062, 33.75388,
    33.44107, 32.36649, 31.65404, 31.78377, 32.25427, 32.36439, 32.18393,
    32.62186, 30.61722,
  44.20086, 44.24883, 44.11446, 43.7757, 44.02849, 46.44106, 46.92691,
    41.89116, 38.35082, 38.20736, 37.49605, 36.92612, 36.57606, 36.99971,
    37.71948, 37.57384, 36.23957, 34.48596, 33.49134, 32.25623, 31.48773,
    31.21774, 30.9886, 30.76764, 30.79498, 31.2346, 31.33133, 30.64889,
    29.90536, 29.01773,
  23.93595, 23.97888, 24.01945, 24.06172, 24.03997, 24.04211, 24.0561,
    24.08944, 24.16367, 24.27371, 25.17597, 25.41694, 24.28555, 24.43878,
    24.59, 24.21446, 24.12485, 24.17149, 24.23446, 24.86063, 25.22455,
    24.63281, 24.58371, 25.19865, 25.59002, 25.26635, 27.89647, 29.94059,
    26.18404, 24.75833,
  24.42666, 24.53526, 24.2177, 24.50128, 24.34433, 24.1762, 24.26759,
    24.3645, 24.47357, 24.66146, 25.09063, 25.70012, 26.06984, 25.35875,
    24.91284, 25.02017, 24.44783, 24.55502, 25.09635, 25.64021, 25.57513,
    25.05705, 25.12946, 26.16988, 30.48132, 31.70878, 28.48441, 31.87427,
    26.96148, 25.34797,
  24.38615, 24.39051, 24.32875, 24.37952, 24.33023, 24.32684, 24.37808,
    24.48693, 24.61497, 24.68795, 24.82382, 25.26385, 25.60052, 26.11093,
    26.3177, 25.43416, 25.36927, 25.82946, 25.88842, 26.18351, 27.11454,
    28.52152, 29.57478, 29.4307, 34.37626, 37.58881, 30.86468, 31.19162,
    26.76948, 25.93339,
  24.55236, 24.54145, 24.72994, 24.93071, 25.20104, 25.73866, 25.85872,
    25.62165, 25.66623, 25.92232, 26.06774, 26.43359, 26.35404, 25.98509,
    27.13224, 28.33626, 27.68832, 26.43892, 26.81447, 27.4645, 30.12488,
    31.56745, 30.1422, 34.92587, 37.52503, 33.15289, 33.73985, 30.38071,
    26.83319, 25.2129,
  25.47063, 25.1722, 25.52273, 25.90175, 26.21155, 26.38271, 26.39704,
    26.29539, 26.78069, 27.22907, 27.03877, 27.03957, 27.00302, 27.4487,
    28.37218, 29.08353, 28.30498, 27.35822, 28.0111, 32.88174, 35.08451,
    29.19519, 28.95079, 30.90896, 32.98065, 32.53063, 30.66974, 31.04736,
    31.84495, 27.12444,
  26.11629, 26.3335, 27.09839, 28.26191, 28.27211, 27.6082, 27.69491,
    27.59042, 27.22071, 27.35203, 27.64729, 29.52502, 31.96885, 32.23314,
    32.03331, 39.33921, 47.51958, 37.8569, 31.29752, 33.27569, 31.44406,
    27.68046, 28.11593, 29.07544, 31.80371, 31.5278, 33.92306, 47.91169,
    43.75671, 26.41155,
  27.3222, 27.81151, 28.66401, 29.736, 30.01799, 29.92244, 30.82288,
    32.55219, 32.90215, 32.95946, 33.61802, 33.13837, 31.87097, 32.10433,
    37.79322, 45.88966, 42.34405, 33.76562, 30.73252, 30.42035, 28.79554,
    27.63739, 28.09554, 30.40011, 32.08347, 29.67935, 39.42991, 57.14645,
    43.90355, 24.73222,
  28.87652, 29.57966, 30.78433, 32.10669, 32.31435, 34.60932, 37.26999,
    35.1046, 33.27343, 33.29575, 32.84813, 31.59321, 30.20221, 30.26431,
    32.18042, 33.9626, 32.77569, 31.24352, 29.10131, 28.65223, 27.95299,
    27.55048, 28.78052, 31.12571, 31.04144, 29.42305, 42.18932, 49.59116,
    31.72896, 25.12896,
  32.48838, 33.18386, 34.52536, 35.18373, 35.59515, 37.56968, 36.58372,
    34.60798, 34.33767, 33.93383, 32.73011, 31.17759, 30.22955, 33.57298,
    36.26611, 32.20039, 31.52103, 33.15956, 33.10032, 30.38492, 27.95873,
    29.54683, 33.82118, 34.82984, 31.04486, 31.55702, 37.86627, 36.82811,
    27.2305, 25.10335,
  37.8236, 40.32884, 41.92398, 43.50019, 42.87978, 39.0727, 34.51604,
    34.24559, 33.37238, 32.79191, 33.52304, 37.11721, 38.47828, 37.0215,
    34.58736, 34.61673, 35.26807, 35.66712, 34.12244, 32.11469, 32.17397,
    32.85417, 33.78772, 31.88137, 37.78571, 49.43658, 41.14878, 28.35417,
    25.55545, 24.18582,
  53.68745, 56.33025, 51.05632, 44.95489, 43.21722, 42.19865, 38.35971,
    40.18382, 42.04391, 49.3956, 54.7189, 38.30866, 33.40251, 32.41696,
    31.66535, 32.40529, 33.45906, 33.27894, 32.23109, 31.98338, 34.4825,
    33.88991, 30.85018, 28.65149, 32.61715, 36.69208, 30.67978, 25.07413,
    24.63458, 24.0155,
  70.1658, 55.6482, 58.52454, 60.52929, 58.87302, 50.90567, 53.34104,
    49.97244, 42.04243, 45.74048, 45.20199, 31.84435, 32.87452, 33.80984,
    31.3124, 31.73892, 30.97088, 30.75804, 30.45403, 30.90504, 33.68725,
    32.51696, 28.08207, 31.57308, 33.9515, 27.26908, 24.5852, 24.92578,
    24.8327, 24.24279,
  79.86061, 75.69415, 91.80194, 94.53925, 96.77799, 85.21648, 65.16806,
    44.57215, 43.60009, 40.3343, 37.6506, 31.3414, 35.73614, 38.00792,
    32.8861, 31.83679, 31.4154, 30.83829, 30.02081, 32.08635, 33.6893,
    30.43366, 27.57896, 32.31216, 34.13981, 26.21479, 24.78948, 25.08971,
    25.38604, 24.60284,
  84.88773, 96.06633, 97.221, 96.5209, 82.49846, 71.94476, 69.78194,
    65.42428, 56.0365, 50.87997, 58.79637, 57.75335, 59.26022, 57.65083,
    50.3703, 39.46783, 32.14725, 33.79354, 34.91462, 35.71381, 32.86679,
    31.6572, 33.70163, 29.63826, 27.08115, 25.44223, 24.82677, 24.61659,
    25.04358, 24.56336,
  63.12213, 67.7029, 63.15683, 58.73817, 52.27504, 59.53455, 83.75964,
    81.16848, 71.87535, 72.00959, 69.05421, 53.97736, 42.68287, 47.96225,
    50.74763, 36.20512, 36.28902, 36.21544, 39.38689, 40.73112, 36.05102,
    32.35333, 28.8204, 26.22986, 25.15775, 25.50838, 24.93398, 24.54308,
    24.49697, 24.22904,
  50.03897, 48.09119, 46.60352, 44.76535, 44.82082, 50.28234, 57.36984,
    55.68978, 52.84107, 50.6543, 46.88291, 39.30793, 34.65606, 38.2303,
    38.15989, 35.39324, 36.91464, 35.19736, 36.44457, 36.36592, 30.32301,
    27.47747, 25.42261, 25.36481, 25.68827, 25.46762, 25.01017, 24.64422,
    24.43067, 24.14745,
  45.2494, 42.95397, 41.81485, 41.6814, 43.01822, 44.2271, 44.65151,
    44.45732, 42.85242, 40.64686, 36.29158, 35.48716, 39.61817, 38.1038,
    35.54029, 35.63507, 34.85135, 32.75659, 34.67949, 33.90241, 26.32324,
    26.25219, 25.8997, 25.53008, 25.41678, 25.45702, 24.95076, 24.37192,
    24.30679, 24.13134,
  40.73288, 40.35611, 40.05767, 40.75938, 41.09626, 41.61843, 41.43708,
    40.65067, 39.60547, 36.46161, 35.73638, 38.4674, 38.89534, 38.32445,
    39.75944, 37.22385, 32.50471, 29.74453, 32.75701, 32.04676, 26.39132,
    26.66807, 26.38979, 25.89383, 25.01164, 25.04251, 24.78469, 24.18385,
    24.11937, 24.03561,
  41.4442, 41.66648, 40.23372, 39.3065, 39.1117, 38.55347, 38.0335, 37.50502,
    36.16093, 34.55296, 36.59243, 36.96357, 32.67855, 33.30416, 34.32462,
    33.07037, 32.56162, 32.78339, 35.71718, 35.34137, 30.21286, 27.85695,
    26.70112, 26.08178, 24.9187, 24.6805, 24.54681, 24.1866, 24.07467,
    24.00002,
  42.05592, 41.58794, 39.61634, 37.66307, 37.15327, 36.63596, 36.18028,
    35.63953, 34.7723, 36.10858, 36.96805, 32.57826, 29.93125, 30.01743,
    29.86725, 29.14738, 30.50791, 32.67411, 35.03456, 36.01731, 33.37012,
    29.79362, 26.96443, 26.20409, 25.28019, 24.71084, 24.4789, 24.22348,
    24.08561, 24.00998,
  40.96018, 40.2787, 38.26322, 36.49652, 35.8842, 35.67252, 35.35896,
    34.79764, 34.63811, 35.83821, 33.52829, 28.90308, 29.03599, 29.34404,
    29.06975, 28.3912, 28.72017, 29.51589, 31.01377, 31.60229, 31.07265,
    30.42627, 28.69845, 26.82894, 25.63537, 24.99978, 24.49526, 24.23181,
    24.10343, 24.01209,
  40.88793, 39.04874, 37.37037, 36.23269, 35.77596, 35.02465, 34.66544,
    33.88631, 34.46187, 34.2632, 30.16885, 27.52488, 28.32177, 28.56538,
    28.39627, 28.20704, 27.89254, 27.8196, 28.01136, 27.73979, 28.94688,
    29.81261, 29.50412, 29.96746, 28.06491, 25.71859, 24.64925, 24.40607,
    24.15459, 24.02926,
  39.83947, 38.48507, 36.62408, 35.55003, 36.02804, 36.09279, 35.21697,
    33.66409, 33.86481, 32.28238, 28.17933, 27.30938, 27.86371, 28.11552,
    27.82405, 28.21349, 28.16834, 27.14857, 26.56848, 26.41747, 27.87378,
    28.43453, 27.57315, 29.31464, 29.55551, 26.83667, 24.92967, 24.89299,
    24.47818, 24.07171,
  39.0805, 37.87144, 37.09905, 36.66056, 36.61785, 36.35016, 36.44463,
    35.99617, 36.24766, 32.54459, 27.94429, 28.06203, 28.60925, 29.06171,
    28.91784, 28.96685, 29.13942, 28.23051, 26.85346, 26.67807, 27.22426,
    27.2256, 26.78653, 27.16962, 28.33096, 28.42267, 26.60882, 25.31149,
    24.87962, 24.24653,
  38.56907, 38.74812, 36.47601, 35.75674, 36.18083, 36.16737, 35.65507,
    35.5655, 36.76672, 33.17269, 28.27392, 28.57299, 29.14147, 29.38046,
    29.31443, 29.46294, 29.27107, 29.05044, 27.81647, 26.55093, 26.94306,
    27.33739, 27.09838, 26.32245, 25.94182, 27.27322, 27.51011, 26.19803,
    25.77184, 24.74037,
  38.58078, 40.14955, 39.45848, 37.58601, 36.38503, 35.54445, 36.5239,
    37.55704, 35.80673, 31.96357, 29.07247, 29.27159, 29.94228, 29.43055,
    28.76357, 28.8215, 28.82809, 29.00084, 28.20447, 26.83609, 27.31536,
    27.67382, 26.59566, 25.68472, 25.50093, 26.19248, 27.60222, 26.88121,
    25.64441, 24.65831,
  39.6483, 41.13264, 38.46962, 36.74921, 35.99246, 35.00822, 36.4639,
    37.00968, 33.64015, 30.20469, 29.25978, 29.46577, 29.71336, 29.04745,
    28.51337, 28.36198, 28.29173, 28.58003, 27.94656, 26.68758, 27.51518,
    29.2292, 29.32299, 27.8942, 27.21957, 27.44035, 29.16726, 28.93862,
    25.75266, 24.09175,
  39.22126, 39.48335, 37.54692, 36.90427, 37.19152, 36.5595, 37.16772,
    35.61414, 31.23733, 29.56285, 28.87426, 29.06659, 29.22756, 28.85716,
    29.00826, 28.70086, 28.06878, 28.19999, 28.2857, 28.13006, 29.75036,
    30.67757, 29.60313, 28.26247, 27.75127, 28.0103, 28.50383, 30.40268,
    28.76715, 24.90212,
  36.69425, 35.8364, 36.4096, 37.74844, 38.63166, 39.75803, 38.38764,
    34.09872, 30.76728, 29.66601, 28.05832, 27.39125, 27.36743, 27.91959,
    29.06137, 29.6147, 29.75557, 30.15017, 29.18228, 27.94403, 28.28695,
    27.97217, 26.93225, 26.30316, 26.53847, 27.11479, 27.2777, 27.2898,
    27.76793, 25.57898,
  35.77115, 35.9079, 35.93686, 35.88625, 36.39382, 39.14098, 39.67759,
    34.41795, 30.62747, 30.19626, 29.74582, 29.77032, 29.89953, 30.59632,
    31.45391, 31.47092, 30.29909, 28.74926, 27.75504, 26.62007, 25.9906,
    25.76781, 25.60087, 25.4994, 25.62494, 26.16861, 26.3433, 25.75066,
    25.17173, 24.31779,
  17.53905, 17.56769, 17.59841, 17.62405, 17.60214, 17.60248, 17.61409,
    17.63196, 17.67151, 17.73347, 18.5144, 18.68992, 17.79941, 17.94105,
    18.05134, 17.73207, 17.65159, 17.68362, 17.69771, 18.19504, 18.509,
    18.04187, 17.95347, 18.41139, 18.6891, 18.35112, 20.59023, 22.32188,
    19.47744, 18.23151,
  17.86466, 17.92827, 17.70559, 17.93772, 17.80659, 17.66288, 17.72053,
    17.77913, 17.85851, 18.00771, 18.39124, 18.93103, 19.22836, 18.63131,
    18.29216, 18.31816, 17.83109, 17.88605, 18.29201, 18.72598, 18.69197,
    18.19483, 18.16979, 18.91154, 22.67556, 23.52663, 21.44389, 24.74181,
    20.43818, 18.86494,
  17.80673, 17.81281, 17.75657, 17.80491, 17.76366, 17.7345, 17.75803,
    17.83239, 17.92567, 17.99402, 18.10821, 18.50867, 18.7909, 19.19063,
    19.3128, 18.51772, 18.41114, 18.76154, 18.74198, 18.88939, 19.55793,
    20.71378, 21.68401, 21.35558, 26.12255, 29.25916, 23.92796, 24.39831,
    20.31127, 19.40691,
  17.83557, 17.82956, 17.96958, 18.10901, 18.32758, 18.74862, 18.80025,
    18.57754, 18.61571, 18.85639, 18.99566, 19.33678, 19.20313, 18.84346,
    19.72016, 20.61066, 19.99907, 18.93584, 19.08257, 19.42248, 21.69647,
    23.13112, 22.14804, 26.4847, 28.71391, 25.80869, 27.02537, 23.84174,
    20.2314, 18.71771,
  18.33529, 18.05447, 18.30706, 18.59972, 18.86727, 19.01844, 19.00019,
    18.86746, 19.3031, 19.71256, 19.6311, 19.59923, 19.42558, 19.67485,
    20.36978, 20.81403, 19.9736, 19.23673, 19.69188, 24.39436, 26.46267,
    21.33536, 21.2174, 23.19105, 24.87844, 24.6829, 23.90164, 24.15536,
    24.73685, 20.42011,
  18.39658, 18.47979, 19.14703, 20.14985, 20.14057, 19.57064, 19.6188,
    19.45068, 19.11606, 19.21804, 19.3443, 20.97044, 23.02255, 23.20838,
    22.72267, 29.26721, 36.4876, 28.33219, 22.81875, 25.11473, 23.62952,
    20.09157, 20.50554, 21.20143, 23.64453, 23.65456, 26.02302, 38.08067,
    34.51887, 19.74598,
  18.85134, 19.19352, 19.95831, 20.88808, 21.02713, 20.68926, 21.29427,
    22.74249, 23.01909, 23.03342, 23.69842, 23.52176, 22.66912, 22.75613,
    27.56139, 35.17736, 33.16513, 25.32699, 22.74831, 22.53531, 21.01974,
    20.00556, 20.46871, 22.69573, 24.3047, 22.15342, 31.56818, 47.5556,
    35.19535, 18.19095,
  19.69568, 20.08767, 20.99367, 21.9837, 21.9997, 23.92743, 26.1704, 24.3135,
    22.84847, 23.02571, 22.95536, 22.13016, 21.19263, 21.41736, 23.52781,
    25.48636, 24.40037, 22.89599, 21.2584, 20.95802, 20.39229, 19.99251,
    21.20018, 23.56534, 23.55527, 22.01956, 34.91738, 41.7446, 24.83789,
    18.50998,
  22.22626, 22.51936, 23.58323, 24.04815, 24.44428, 26.36148, 25.65176,
    23.84831, 23.7189, 23.62901, 22.88752, 21.82174, 21.1676, 24.20001,
    26.4922, 23.30185, 23.11342, 24.85358, 24.76282, 22.38281, 20.24698,
    21.62476, 25.62132, 26.61615, 23.28212, 23.71437, 30.46828, 29.67908,
    20.56695, 18.58808,
  26.18888, 27.98099, 29.39425, 30.6541, 30.58439, 27.87062, 24.24651,
    23.88686, 23.21012, 22.43786, 23.11922, 26.42082, 28.11516, 27.72413,
    26.01854, 25.99685, 26.76786, 27.34311, 25.94275, 24.12182, 23.95648,
    24.72561, 25.96439, 24.50755, 29.64656, 39.86073, 33.11665, 21.6827,
    19.09294, 17.79994,
  38.07267, 41.13609, 37.60334, 33.16462, 31.99846, 30.83582, 27.25821,
    28.60372, 29.91014, 36.37714, 40.76192, 28.1738, 24.70839, 24.18882,
    23.46666, 24.26349, 25.44755, 25.3767, 24.36659, 24.06737, 26.42003,
    26.25835, 23.39496, 21.40214, 25.66284, 30.15829, 24.41123, 18.60738,
    18.16625, 17.61567,
  52.68788, 41.62014, 43.64461, 45.10575, 43.49272, 37.55333, 40.3605,
    37.58959, 31.11124, 35.28221, 35.33755, 22.89561, 23.91406, 24.8577,
    23.07349, 23.49393, 22.94277, 22.89349, 22.58302, 23.25486, 26.15993,
    25.15843, 21.00145, 24.17941, 26.44147, 20.70527, 18.1294, 18.434,
    18.38372, 17.83483,
  60.76628, 56.46551, 74.45927, 78.94647, 77.29792, 67.63586, 52.22373,
    35.45057, 33.02414, 31.14731, 28.41387, 21.33488, 25.92755, 28.62187,
    24.26112, 23.51565, 23.52979, 22.92975, 22.37984, 24.76505, 26.63788,
    23.45445, 20.67931, 25.6232, 27.44246, 19.77175, 18.29574, 18.62016,
    18.94022, 18.17733,
  66.80432, 93.90952, 92.67827, 86.67216, 73.75799, 63.56599, 57.19762,
    51.63227, 43.43272, 37.90723, 43.94244, 43.00064, 45.91217, 45.21048,
    38.76371, 30.5294, 24.22533, 25.84974, 27.17773, 28.20803, 25.87494,
    24.73903, 26.655, 23.41683, 20.79701, 18.88085, 18.37803, 18.21594,
    18.6574, 18.15571,
  50.23586, 58.069, 55.59561, 52.3893, 45.69044, 49.02496, 67.44071,
    65.78884, 56.17658, 56.32103, 55.44242, 43.04053, 33.38841, 38.54736,
    40.96205, 28.34189, 27.88263, 28.15262, 30.82541, 32.1584, 28.90404,
    25.83448, 22.80981, 19.96336, 18.48929, 18.88799, 18.46222, 18.11401,
    18.10964, 17.84166,
  39.67821, 39.17572, 38.35191, 36.53461, 35.51985, 39.72826, 46.52975,
    44.82819, 41.7014, 40.73745, 38.2614, 30.32431, 25.43019, 29.49355,
    29.71371, 27.04988, 28.86409, 27.513, 28.57714, 28.72051, 23.99932,
    21.2846, 18.99666, 18.8199, 19.07008, 18.86777, 18.52048, 18.21331,
    18.02895, 17.75484,
  37.01578, 35.38762, 33.78209, 32.90497, 33.47651, 34.57947, 35.05532,
    34.72582, 33.45479, 31.52235, 27.30248, 26.40518, 29.82778, 28.42862,
    27.11563, 27.48389, 27.19345, 25.41817, 26.79101, 25.99058, 19.81441,
    19.63813, 19.39251, 19.0834, 18.9088, 18.90807, 18.46253, 17.9725,
    17.91717, 17.73935,
  33.03484, 32.01809, 31.04284, 31.46804, 31.95389, 32.78738, 33.04217,
    32.50863, 31.29608, 27.82301, 26.69942, 29.49863, 30.10484, 29.57445,
    31.09812, 29.47095, 25.54511, 22.97132, 25.37504, 24.47615, 19.62112,
    19.93401, 19.8294, 19.42812, 18.5488, 18.56759, 18.31421, 17.7807,
    17.74605, 17.65097,
  32.46492, 32.31206, 30.99876, 30.50023, 30.77253, 30.75194, 30.55031,
    29.8598, 28.07403, 26.12401, 28.19278, 28.98213, 25.40251, 26.13834,
    27.12418, 26.07101, 25.50145, 25.5277, 27.53188, 26.63721, 22.70057,
    21.04012, 20.11443, 19.56309, 18.44232, 18.23075, 18.10452, 17.77893,
    17.70522, 17.62498,
  32.85429, 32.70944, 31.13232, 29.66474, 29.59279, 29.31315, 28.88424,
    28.14274, 27.073, 28.27393, 29.44332, 25.76616, 23.18151, 23.23294,
    22.98799, 22.25864, 23.46684, 25.44422, 26.97714, 27.47441, 25.8479,
    22.99084, 20.32805, 19.64062, 18.79471, 18.26081, 18.06192, 17.81623,
    17.70643, 17.63507,
  32.41764, 32.3462, 30.56538, 29.07021, 28.70261, 28.59329, 28.36098,
    27.89671, 27.79985, 29.16441, 27.30593, 22.68942, 22.41251, 22.36177,
    21.82331, 21.19467, 21.57421, 22.48139, 23.64149, 24.13909, 24.1805,
    23.74034, 21.97713, 20.22683, 19.10178, 18.50405, 18.06656, 17.82232,
    17.71332, 17.63249,
  32.92094, 31.71447, 30.09504, 29.10118, 28.85017, 28.44805, 28.49716,
    28.13741, 28.66134, 28.41014, 24.35522, 21.17265, 21.48318, 21.45423,
    21.15756, 21.08006, 20.90523, 20.87326, 21.20448, 21.11655, 22.2629,
    22.81118, 22.09175, 22.46723, 21.02902, 19.05965, 18.18856, 17.9379,
    17.731, 17.63409,
  32.50748, 31.49718, 29.7454, 28.90395, 29.65312, 30.14265, 29.88805,
    28.68211, 28.59977, 26.66381, 22.1906, 20.67328, 20.8409, 20.95495,
    20.73025, 21.20936, 21.19364, 20.27547, 19.88528, 19.81436, 21.17894,
    21.42459, 20.30184, 22.03014, 22.3781, 19.94778, 18.4263, 18.3849,
    18.01917, 17.66542,
  32.02919, 31.20404, 30.5048, 30.46979, 31.0018, 31.22266, 31.41195,
    30.6408, 30.16518, 26.28774, 21.60809, 21.18762, 21.54082, 21.94863,
    21.84065, 21.92394, 21.97618, 21.03266, 19.96704, 19.95493, 20.43183,
    20.30984, 19.79197, 20.22096, 21.28881, 21.35115, 19.91282, 18.79189,
    18.40688, 17.82192,
  32.12574, 32.9334, 30.84374, 30.3342, 30.95358, 30.95244, 30.38929,
    29.90061, 30.50291, 26.77118, 21.85768, 21.72338, 22.07461, 22.37169,
    22.37682, 22.38626, 21.94833, 21.52094, 20.66254, 19.86929, 20.08258,
    20.28763, 20.13696, 19.50067, 19.29083, 20.52163, 20.75369, 19.55107,
    19.2107, 18.25474,
  32.72162, 34.89743, 33.57644, 31.85027, 30.80677, 29.93447, 30.49336,
    31.28363, 29.74831, 25.85599, 22.66767, 22.39932, 22.78536, 22.42615,
    21.81334, 21.76941, 21.51191, 21.45527, 21.04302, 20.15877, 20.39963,
    20.58729, 19.73248, 18.98259, 18.85732, 19.47158, 20.76839, 20.13436,
    19.16114, 18.1995,
  33.78154, 35.66697, 33.04199, 31.11606, 30.19523, 29.18578, 30.54621,
    31.13373, 28.03684, 24.44694, 23.0206, 22.64883, 22.60216, 22.034,
    21.48886, 21.3354, 21.13684, 21.22435, 20.90721, 20.05262, 20.46175,
    21.65109, 21.67652, 20.69456, 20.40599, 20.58154, 22.27217, 21.9948,
    19.15769, 17.70642,
  33.37934, 33.86808, 31.64605, 30.71979, 30.98028, 30.40159, 31.11936,
    29.85094, 25.97232, 23.85807, 22.64474, 22.20241, 21.99701, 21.73826,
    21.9104, 21.65216, 20.99372, 20.92592, 21.18268, 21.27344, 22.21177,
    22.67126, 21.97094, 21.12738, 20.99095, 21.17531, 21.72391, 23.38463,
    21.72985, 18.34132,
  30.71314, 29.83063, 30.19233, 31.54573, 32.51169, 33.35557, 32.27351,
    28.55442, 25.37876, 23.81421, 21.79396, 20.70297, 20.4939, 20.82925,
    21.58472, 21.88634, 21.90442, 22.25287, 21.78866, 21.12149, 21.34882,
    21.06426, 20.17133, 19.67242, 19.9361, 20.40676, 20.51011, 20.62262,
    21.11629, 18.97288,
  29.35081, 29.44375, 29.7642, 30.14917, 30.63655, 32.87382, 33.18591,
    28.52113, 24.89185, 23.85592, 22.80204, 22.41323, 22.48033, 22.73591,
    23.06901, 23.1973, 22.3859, 21.31716, 20.67563, 19.8906, 19.40033,
    19.25407, 19.10171, 19.001, 19.11893, 19.60346, 19.71061, 19.13783,
    18.71213, 17.93273,
  14.11567, 14.14084, 14.16363, 14.17743, 14.17231, 14.16359, 14.16312,
    14.18436, 14.22468, 14.25901, 14.96458, 15.07712, 14.31429, 14.48363,
    14.58057, 14.28841, 14.22436, 14.2373, 14.2371, 14.69902, 14.94822,
    14.52286, 14.44185, 14.84281, 15.00108, 14.65065, 16.7939, 18.26198,
    15.89233, 14.73157,
  14.42409, 14.45083, 14.25383, 14.46946, 14.35248, 14.21124, 14.24362,
    14.28616, 14.34532, 14.48566, 14.87887, 15.35456, 15.58653, 15.06612,
    14.80146, 14.77915, 14.35321, 14.39389, 14.7621, 15.19471, 15.12434,
    14.5487, 14.4705, 15.08815, 18.43641, 18.97504, 17.77026, 20.64552,
    16.81593, 15.31498,
  14.38479, 14.38719, 14.31085, 14.3588, 14.30149, 14.24206, 14.25453,
    14.30841, 14.40133, 14.46051, 14.54754, 14.94204, 15.23753, 15.58994,
    15.62409, 14.89779, 14.79589, 15.09135, 15.06393, 15.12152, 15.5847,
    16.56017, 17.40771, 16.93373, 21.43373, 24.21312, 19.78561, 20.31558,
    16.65218, 15.82655,
  14.34591, 14.32439, 14.46652, 14.59105, 14.78661, 15.18263, 15.21603,
    14.95065, 14.9448, 15.1596, 15.27517, 15.6043, 15.41803, 15.14942,
    15.9294, 16.66343, 16.027, 15.02845, 15.01956, 15.13585, 17.23353,
    18.57641, 17.79641, 21.46019, 23.30475, 21.42436, 22.60346, 19.89358,
    16.52735, 15.19964,
  14.70888, 14.44929, 14.67746, 14.95884, 15.24031, 15.39751, 15.32201,
    15.11863, 15.56611, 16.0464, 16.01665, 15.82202, 15.48064, 15.65044,
    16.25574, 16.57677, 15.55284, 14.79214, 15.15729, 19.39916, 21.1298,
    17.00058, 16.93953, 18.89732, 20.43864, 20.22188, 19.67374, 20.11279,
    20.42464, 16.49252,
  14.62413, 14.63326, 15.32251, 16.35209, 16.39217, 15.84538, 15.71938,
    15.46369, 15.20995, 15.31694, 15.31123, 16.70101, 18.35553, 18.4931,
    17.78219, 23.50486, 29.36851, 22.34091, 17.94586, 20.44423, 19.1482,
    15.87348, 16.37738, 17.03166, 19.29411, 19.02427, 21.0738, 32.14194,
    29.31452, 16.04962,
  14.69902, 15.01065, 15.83741, 16.84206, 17.06964, 16.5939, 16.89694,
    18.23709, 18.46233, 18.3462, 18.97156, 18.77522, 17.92196, 17.78399,
    22.40944, 29.66195, 27.77722, 20.41727, 18.22212, 18.20247, 16.80914,
    15.89484, 16.27079, 18.10143, 19.53114, 17.46937, 25.9306, 40.87666,
    30.45693, 14.69576,
  14.8804, 15.22505, 16.15946, 17.08772, 17.02081, 18.83804, 20.78477,
    19.00896, 17.78417, 17.96216, 18.02995, 17.22244, 16.2717, 16.41878,
    18.95876, 21.13605, 19.826, 18.30031, 16.99945, 16.76427, 16.24499,
    15.89021, 16.81887, 18.8084, 18.86067, 17.18849, 29.49571, 36.26391,
    20.8579, 14.90866,
  16.27941, 16.44261, 17.50119, 17.76221, 18.14664, 20.29595, 19.66376,
    17.74289, 17.80466, 17.99839, 17.489, 16.6298, 16.19073, 19.18714,
    21.22755, 18.54844, 18.41134, 19.84835, 19.7412, 17.71822, 15.92848,
    16.99974, 20.39745, 21.34284, 18.59347, 18.60812, 25.14662, 24.93894,
    16.64189, 15.03312,
  18.38377, 19.74044, 21.25106, 22.45423, 22.63849, 20.27835, 17.16795,
    16.94406, 16.72891, 16.28219, 17.28236, 20.57083, 22.18581, 22.0812,
    21.11544, 21.0876, 21.67879, 22.15403, 21.2639, 19.91228, 19.61755,
    20.45365, 21.7479, 20.4104, 24.65729, 33.58508, 28.10026, 17.99651,
    15.60694, 14.38284,
  27.06738, 29.86495, 27.43008, 23.5637, 22.99221, 22.29673, 19.38041,
    20.86478, 22.42107, 28.48461, 32.03782, 22.39332, 19.89405, 19.54299,
    19.03152, 19.95392, 21.20536, 21.2426, 20.41823, 20.29521, 22.52102,
    22.44767, 19.78542, 17.77431, 21.90197, 26.63099, 21.26206, 15.27484,
    14.72163, 14.18663,
  39.01203, 29.65272, 31.14324, 32.34411, 31.22775, 27.41812, 30.4488,
    28.57798, 23.63688, 28.44053, 28.67652, 18.17913, 19.19469, 20.37623,
    19.13628, 19.57321, 19.14749, 19.21219, 19.00844, 19.695, 22.58857,
    21.59372, 17.44302, 20.38597, 22.74257, 17.46892, 14.73577, 14.91496,
    14.92112, 14.40821,
  44.17113, 40.60612, 57.73481, 62.5946, 62.22275, 54.00368, 40.64814,
    27.06619, 25.52522, 24.78332, 22.11356, 16.58329, 21.34585, 24.06283,
    20.38157, 19.70457, 19.74811, 19.18939, 18.68135, 21.24531, 23.26847,
    20.01842, 17.15759, 22.12264, 24.09951, 16.36674, 14.76936, 15.11479,
    15.45069, 14.73697,
  52.5913, 76.69294, 77.45304, 71.51892, 60.30114, 51.80733, 46.46904,
    40.72626, 33.90545, 30.47345, 36.06732, 35.67098, 38.93446, 38.92915,
    33.52645, 25.8622, 20.23241, 21.69119, 23.0117, 24.27135, 22.31532,
    21.14884, 23.091, 20.24122, 17.60258, 15.36411, 14.87284, 14.76027,
    15.21755, 14.73555,
  39.51302, 47.94828, 45.99981, 42.82278, 36.53428, 40.42467, 56.85472,
    55.34956, 46.52109, 47.43432, 47.90057, 36.98975, 28.63403, 33.64162,
    36.02121, 24.15427, 23.34513, 23.54171, 25.4722, 26.9923, 24.96163,
    22.27073, 19.85108, 16.78289, 14.95918, 15.39437, 15.00264, 14.66563,
    14.68347, 14.43682,
  29.30118, 29.35657, 29.16125, 28.10337, 27.3642, 32.21083, 39.65732,
    37.71338, 35.15003, 35.54005, 33.09888, 25.77643, 21.17681, 25.43795,
    25.62196, 22.68313, 24.44422, 23.0191, 23.4395, 23.87622, 20.51744,
    18.10661, 15.68326, 15.45685, 15.63922, 15.39338, 15.03848, 14.77391,
    14.61136, 14.33727,
  27.37795, 26.49769, 25.36245, 24.65569, 25.17589, 26.40532, 27.32405,
    27.09899, 26.65289, 25.84024, 22.26196, 22.13885, 25.06093, 23.58141,
    22.88736, 23.1473, 23.13426, 21.24324, 21.88302, 21.34844, 16.3491,
    16.25034, 15.95782, 15.72224, 15.5106, 15.42148, 14.99638, 14.54759,
    14.50049, 14.32904,
  24.57916, 23.80849, 22.81678, 23.11327, 23.68317, 24.72274, 25.4647,
    25.5736, 25.05674, 22.6796, 21.93287, 25.02993, 25.98696, 25.14926,
    26.72928, 25.32469, 21.75392, 19.20751, 21.04495, 20.21207, 16.03142,
    16.32142, 16.19313, 15.90485, 15.14097, 15.10535, 14.88173, 14.36755,
    14.33332, 14.23935,
  24.20417, 24.0297, 22.74596, 22.42085, 22.93605, 23.34567, 23.67814,
    23.56522, 22.47095, 21.19356, 23.43122, 24.75344, 21.82452, 22.52604,
    23.49252, 22.42272, 21.65309, 21.45337, 22.85043, 21.61352, 18.38596,
    17.15175, 16.34219, 15.94728, 14.97888, 14.77374, 14.67992, 14.3566,
    14.28379, 14.20802,
  24.56468, 24.50824, 23.16499, 22.05348, 22.29772, 22.32509, 22.25674,
    22.00123, 21.42681, 22.88321, 24.54162, 21.86495, 19.71612, 19.81303,
    19.51794, 18.83881, 19.81067, 21.48618, 22.28325, 22.24361, 21.18453,
    18.95222, 16.46249, 15.97396, 15.28347, 14.78941, 14.61479, 14.38707,
    14.27692, 14.21019,
  24.20773, 24.46031, 23.11348, 21.93451, 21.79746, 21.79109, 21.71735,
    21.63685, 22.01254, 23.94784, 23.11014, 19.29211, 19.26953, 19.09063,
    18.22271, 17.53373, 17.81447, 18.62784, 19.28375, 19.52587, 20.02812,
    19.8358, 17.92525, 16.52701, 15.66314, 15.06651, 14.62161, 14.38956,
    14.28608, 14.21175,
  24.86122, 24.31, 22.99715, 22.19963, 21.98383, 21.55637, 21.7573, 21.84833,
    22.96034, 23.85474, 20.98106, 17.97388, 18.26433, 18.01396, 17.44548,
    17.26979, 17.10153, 17.03819, 17.3887, 17.44993, 18.54878, 18.90141,
    17.85889, 18.28661, 17.1262, 15.44577, 14.72532, 14.47671, 14.29077,
    14.21026,
  25.00381, 24.45812, 22.81334, 22.02542, 22.60751, 22.99963, 23.15296,
    22.60446, 23.20572, 22.61357, 19.08479, 17.41627, 17.38698, 17.26765,
    16.91971, 17.37187, 17.39392, 16.58804, 16.37602, 16.37271, 17.60097,
    17.66213, 16.30941, 17.96098, 18.322, 16.20267, 14.92288, 14.89142,
    14.55955, 14.24271,
  24.80331, 24.26837, 23.43767, 23.37792, 23.97563, 24.3006, 24.99088,
    24.88518, 24.86403, 22.03557, 18.23626, 17.71502, 17.83057, 18.00634,
    17.79828, 17.98274, 18.05725, 17.17237, 16.34819, 16.4048, 16.74231,
    16.52894, 16.00995, 16.4317, 17.37938, 17.51297, 16.3054, 15.30306,
    14.94918, 14.38208,
  25.03391, 25.71617, 23.814, 23.47061, 24.32863, 24.59855, 24.39361,
    24.14912, 24.95851, 22.25845, 18.22984, 18.05339, 18.18495, 18.38103,
    18.36789, 18.37542, 17.96248, 17.55113, 16.91537, 16.41033, 16.36776,
    16.37243, 16.35133, 15.8914, 15.80836, 17.05331, 17.31535, 16.118,
    15.74778, 14.81487,
  25.64857, 27.93227, 26.60496, 25.03983, 24.49837, 23.83492, 24.17126,
    24.86871, 24.02089, 21.33724, 18.85842, 18.57994, 18.71328, 18.44064,
    17.89952, 17.82243, 17.53224, 17.4606, 17.29727, 16.69181, 16.64117,
    16.69068, 16.04938, 15.46416, 15.42964, 16.12006, 17.46737, 16.78946,
    15.77196, 14.80633,
  26.95615, 29.42636, 26.97349, 24.87167, 23.98442, 22.86453, 24.17535,
    24.89515, 22.50398, 19.97285, 19.28019, 18.9873, 18.75445, 18.22478,
    17.60083, 17.38115, 17.18955, 17.26743, 17.15046, 16.55425, 16.68015,
    17.54771, 17.63311, 17.04951, 17.00559, 17.24691, 19.03123, 18.62941,
    15.70506, 14.29626,
  27.16632, 28.24852, 25.62049, 24.19077, 24.33098, 23.51589, 24.21762,
    23.56422, 20.69356, 19.50864, 19.0955, 18.67944, 18.23943, 17.94651,
    17.98489, 17.69538, 17.07933, 16.94111, 17.3378, 17.71132, 18.12976,
    18.26038, 17.91091, 17.5226, 17.72239, 17.89719, 18.47069, 20.00679,
    18.20985, 14.88076,
  25.0578, 23.97824, 23.88619, 25.01545, 25.60148, 25.73851, 24.98425,
    22.29821, 20.13766, 19.57373, 18.27314, 17.28998, 17.00683, 17.1174,
    17.63141, 17.881, 17.82022, 18.09484, 17.9773, 17.64591, 17.70467,
    17.35043, 16.57704, 16.23645, 16.59763, 17.05945, 17.14368, 17.32294,
    17.74142, 15.5412,
  23.53803, 23.22316, 23.46507, 23.95961, 24.25567, 25.74722, 25.85159,
    22.34525, 19.82412, 19.50091, 18.7937, 18.4663, 18.6332, 18.68784,
    18.75361, 18.89432, 18.28977, 17.47649, 17.0518, 16.41713, 15.9526,
    15.85589, 15.66917, 15.57872, 15.71546, 16.18475, 16.30391, 15.72768,
    15.32074, 14.53966,
  12.77768, 12.80534, 12.82791, 12.84049, 12.83763, 12.82756, 12.83013,
    12.84144, 12.87061, 12.88893, 13.5547, 13.62195, 12.91378, 13.08257,
    13.1912, 12.9281, 12.87453, 12.89886, 12.87651, 13.2812, 13.51555,
    13.14769, 13.05953, 13.43574, 13.54418, 13.14987, 15.20195, 16.52934,
    14.45445, 13.40572,
  13.07391, 13.08068, 12.91378, 13.12342, 13.00449, 12.88639, 12.91168,
    12.9348, 12.9782, 13.10441, 13.54201, 13.95964, 14.07628, 13.6096,
    13.43278, 13.38722, 12.99276, 13.0262, 13.36043, 13.81999, 13.79725,
    13.18778, 13.04904, 13.58709, 16.84141, 17.17411, 16.65847, 19.64605,
    15.59646, 14.05747,
  13.07162, 13.07735, 12.99696, 13.06425, 12.97978, 12.89032, 12.89765,
    12.95298, 13.04006, 13.10635, 13.17344, 13.54485, 13.85506, 14.13937,
    14.13574, 13.46002, 13.36404, 13.68543, 13.69496, 13.72822, 14.07463,
    14.87772, 15.73205, 15.1409, 19.85124, 22.62384, 18.58216, 19.32957,
    15.45702, 14.513,
  12.99194, 12.97613, 13.13512, 13.24115, 13.42376, 13.76462, 13.77837,
    13.53419, 13.49288, 13.68357, 13.79117, 14.13643, 13.93656, 13.70492,
    14.3707, 14.9855, 14.49746, 13.64314, 13.53439, 13.48434, 15.53185,
    16.95024, 16.25724, 20.03877, 21.92044, 20.33634, 21.43748, 18.65992,
    15.27032, 13.92241,
  13.30383, 13.07398, 13.29314, 13.57061, 13.86838, 14.06767, 13.96932,
    13.70483, 14.08217, 14.59853, 14.67779, 14.42378, 13.9889, 14.05419,
    14.66638, 15.02975, 13.91915, 13.14107, 13.39105, 17.68641, 19.42744,
    15.61818, 15.45759, 17.85981, 19.36164, 18.80491, 18.51184, 18.63044,
    18.73125, 14.99639,
  13.24437, 13.19151, 13.83502, 14.84304, 14.96104, 14.46371, 14.2985,
    14.00534, 13.78311, 13.92495, 13.81592, 15.07715, 16.59198, 16.74391,
    15.82322, 20.93919, 26.21596, 20.09254, 16.09946, 19.02345, 17.91041,
    14.46605, 15.03818, 15.60135, 17.88169, 17.58406, 19.11183, 29.5894,
    27.37782, 14.75576,
  13.24337, 13.51865, 14.38874, 15.44772, 15.72968, 15.10564, 15.21513,
    16.44838, 16.57315, 16.42072, 17.06425, 17.07582, 16.39464, 16.10316,
    20.40157, 27.77983, 26.50735, 19.08014, 16.82368, 16.82716, 15.44193,
    14.55276, 14.93289, 16.69206, 18.11543, 15.89364, 24.007, 39.16488,
    29.33999, 13.41509,
  13.42053, 13.75356, 14.70221, 15.59512, 15.43025, 17.09055, 18.91579,
    17.33278, 16.27914, 16.45277, 16.62686, 15.73742, 14.61286, 14.58294,
    17.60331, 20.26339, 18.64425, 16.7529, 15.61491, 15.40702, 14.92008,
    14.56654, 15.42575, 17.4244, 17.49796, 15.48838, 28.5605, 35.93834,
    19.96736, 13.54914,
  14.64697, 14.72928, 15.66802, 15.86669, 16.29128, 18.81236, 18.40174,
    16.18215, 16.18307, 16.39604, 15.81589, 14.87118, 14.33075, 17.4988,
    19.59102, 16.98098, 16.9299, 18.34329, 18.18387, 16.27134, 14.55858,
    15.48992, 18.84953, 19.79246, 17.15557, 17.00129, 24.4522, 24.37674,
    15.32477, 13.75548,
  16.48853, 17.58804, 19.08949, 20.3152, 20.75118, 18.61659, 15.64986,
    15.26667, 15.1345, 14.56342, 15.4394, 18.62225, 20.29158, 20.50693,
    19.81524, 19.46404, 19.88405, 20.4986, 19.86876, 18.53614, 18.00521,
    18.96594, 20.51551, 19.21084, 23.06254, 31.73053, 26.80077, 16.97685,
    14.44385, 13.09635,
  23.49836, 26.03094, 24.30065, 21.00455, 20.98004, 20.32848, 17.55155,
    18.99491, 20.07455, 25.47714, 28.85098, 21.075, 18.84671, 18.33451,
    17.55075, 18.51308, 19.80747, 19.88974, 18.97064, 18.83772, 21.06397,
    21.18801, 18.61741, 16.5367, 20.99487, 26.36234, 20.76888, 14.151,
    13.43541, 12.85062,
  34.15771, 25.99588, 27.15652, 28.16005, 27.08377, 23.86093, 26.91494,
    25.69228, 21.55155, 26.60899, 27.16027, 17.03505, 17.62876, 18.70076,
    17.6945, 18.06389, 17.70332, 17.75502, 17.48775, 18.14479, 21.20667,
    20.3615, 16.21299, 19.33138, 21.82201, 16.49084, 13.52374, 13.61866,
    13.6153, 13.0792,
  40.64888, 34.49821, 46.51793, 52.1979, 52.35629, 46.8172, 36.51048,
    24.18484, 23.10888, 22.97504, 20.19925, 14.91138, 19.53156, 22.056,
    18.79371, 18.08546, 18.13778, 17.61134, 17.12772, 19.73181, 21.9129,
    18.8498, 15.86785, 21.60564, 23.77948, 15.34117, 13.48013, 13.8451,
    14.14963, 13.40623,
  47.52148, 67.11755, 70.04116, 69.87425, 65.25032, 55.05478, 40.58976,
    36.51286, 30.09048, 27.62292, 32.84488, 32.73892, 36.68587, 37.05687,
    31.52914, 24.18734, 18.67481, 20.17432, 21.51862, 22.93496, 21.01065,
    20.12775, 22.25105, 19.78983, 16.96543, 14.12722, 13.5702, 13.47344,
    13.93478, 13.41296,
  34.7437, 43.18945, 43.95906, 44.65202, 40.09867, 39.95165, 51.25061,
    51.26881, 42.13866, 43.81762, 45.05554, 35.12806, 27.83825, 32.99804,
    34.70106, 22.85874, 21.87676, 22.04497, 23.89369, 25.67469, 23.90385,
    21.63638, 19.44066, 15.94598, 13.63042, 14.089, 13.66986, 13.34376,
    13.38413, 13.1162,
  24.61398, 25.09677, 26.1612, 25.92221, 24.11609, 28.18629, 36.30676,
    34.09314, 31.88778, 33.62799, 31.79613, 24.37972, 19.67678, 24.26301,
    24.45198, 21.208, 23.14924, 21.68503, 22.03491, 22.89247, 19.9397,
    17.40797, 14.62675, 14.21213, 14.31586, 14.07663, 13.71038, 13.45367,
    13.29533, 13.0102,
  23.30384, 22.91432, 22.16854, 21.20292, 21.17671, 22.36872, 23.4507,
    23.11665, 23.29352, 23.52485, 20.56433, 20.53652, 23.30807, 21.96856,
    21.46009, 21.7655, 22.02272, 20.1146, 20.78812, 20.4429, 15.37724,
    15.1017, 14.74845, 14.47533, 14.24125, 14.10806, 13.64177, 13.22829,
    13.20169, 13.00364,
  21.01666, 20.35814, 19.29056, 19.3915, 19.9406, 21.00805, 21.85669,
    22.28838, 22.05783, 20.22574, 19.61209, 23.08086, 24.78281, 23.95101,
    25.63877, 24.24148, 20.66217, 18.09066, 20.13654, 19.27794, 14.82921,
    14.99135, 14.89028, 14.62847, 13.86623, 13.8406, 13.57218, 13.03023,
    13.01606, 12.9143,
  20.76078, 20.45494, 19.03111, 18.66694, 19.23413, 19.80775, 20.26927,
    20.27853, 19.30549, 18.33918, 21.03288, 23.00522, 20.85205, 21.79848,
    22.92043, 21.74978, 20.65322, 20.10368, 21.56455, 20.37818, 17.07486,
    15.73768, 14.99172, 14.63096, 13.67814, 13.49631, 13.39395, 13.02828,
    12.95273, 12.87197,
  21.15003, 20.96616, 19.51879, 18.38734, 18.70552, 18.75906, 18.71183,
    18.5106, 18.01945, 19.89362, 22.26249, 20.42868, 18.65703, 18.91662,
    18.74117, 18.09432, 18.96383, 20.44998, 21.05736, 21.13108, 20.015,
    17.56691, 15.06529, 14.61812, 13.96674, 13.48293, 13.30083, 13.05265,
    12.94767, 12.8757,
  20.68682, 20.86701, 19.49827, 18.31546, 18.22603, 18.17326, 17.98428,
    17.88144, 18.5793, 21.2828, 21.21068, 18.08995, 18.34893, 18.22946,
    17.33554, 16.56297, 16.71138, 17.43399, 18.06021, 18.50993, 19.14597,
    18.63533, 16.42356, 15.19222, 14.39179, 13.7361, 13.28929, 13.04897,
    12.94538, 12.87394,
  21.2924, 20.68968, 19.3458, 18.53712, 18.24447, 17.73832, 17.86197,
    18.17222, 19.79528, 21.54478, 19.46478, 16.82987, 17.32569, 17.11501,
    16.47914, 16.0986, 15.78839, 15.75659, 16.24587, 16.40807, 17.53328,
    17.71652, 16.59367, 16.84799, 15.63685, 14.05197, 13.36446, 13.1252,
    12.95, 12.8726,
  21.43287, 20.73425, 19.09404, 18.28152, 18.70159, 19.01572, 19.31661,
    19.13814, 20.34958, 20.54868, 17.73422, 16.25084, 16.34801, 16.18937,
    15.75139, 16.10954, 16.09618, 15.35198, 15.21341, 15.21566, 16.46243,
    16.35928, 14.98264, 16.51402, 16.6549, 14.65703, 13.55482, 13.53946,
    13.22844, 12.90871,
  21.11446, 20.48018, 19.5127, 19.38406, 20.02135, 20.47812, 21.5001,
    21.93935, 22.27281, 19.91236, 16.74269, 16.41015, 16.52962, 16.73366,
    16.53672, 16.68492, 16.75376, 15.82305, 15.0174, 15.12806, 15.47835,
    15.14107, 14.53439, 14.92786, 15.80617, 15.93616, 14.83313, 13.9605,
    13.66374, 13.06239,
  21.20318, 21.31889, 19.73667, 19.63712, 20.71083, 21.32071, 21.50134,
    21.57604, 22.46408, 20.04938, 16.50601, 16.60014, 16.90406, 17.18629,
    17.18427, 17.12347, 16.63891, 16.14119, 15.50583, 15.13345, 15.01931,
    14.89716, 14.90458, 14.45668, 14.41549, 15.73178, 15.93556, 14.77562,
    14.50261, 13.48544,
  21.60126, 23.10627, 22.19318, 21.25733, 21.1796, 20.968, 21.3721, 22.02198,
    21.20318, 18.99881, 16.88342, 17.04763, 17.47544, 17.25174, 16.67535,
    16.54784, 16.14567, 16.01137, 15.88165, 15.3262, 15.22423, 15.25804,
    14.66139, 14.10738, 14.07181, 14.76635, 16.16829, 15.46382, 14.5539,
    13.51404,
  22.84555, 24.76395, 23.1578, 21.74501, 20.98419, 20.01016, 21.32972,
    22.03897, 19.64614, 17.54448, 17.33278, 17.56205, 17.54873, 16.9731,
    16.28139, 15.97953, 15.78317, 15.88488, 15.78881, 15.18886, 15.19666,
    16.01439, 16.07255, 15.52645, 15.58553, 15.85743, 17.78378, 17.38794,
    14.45784, 12.99014,
  23.53665, 24.60989, 22.25375, 21.28554, 21.38702, 20.59036, 21.3155,
    20.59696, 17.7954, 17.05454, 17.27994, 17.30869, 16.95666, 16.60836,
    16.61612, 16.25867, 15.67044, 15.59846, 16.03147, 16.3361, 16.57614,
    16.73413, 16.5119, 16.17186, 16.44284, 16.60008, 17.27783, 18.93341,
    16.97503, 13.54186,
  22.05406, 21.12878, 21.10493, 22.38841, 22.76194, 22.64263, 21.97403,
    19.20535, 17.15767, 17.12251, 16.49859, 15.89644, 15.69908, 15.82389,
    16.35939, 16.54601, 16.43962, 16.69627, 16.70097, 16.46482, 16.44896,
    16.09148, 15.31274, 14.97315, 15.37848, 15.89505, 15.96072, 16.22025,
    16.73128, 14.26003,
  21.01201, 20.62247, 21.00944, 21.6701, 21.79604, 22.91406, 22.63411,
    19.09628, 16.92679, 17.03336, 16.7491, 16.71325, 17.00387, 17.25935,
    17.44216, 17.55116, 16.93552, 16.16035, 15.84852, 15.22924, 14.73522,
    14.64508, 14.41674, 14.29386, 14.45569, 15.01708, 15.14937, 14.49279,
    14.16134, 13.27711,
  12.11168, 12.12693, 12.15777, 12.1793, 12.17305, 12.16707, 12.16503,
    12.17672, 12.19864, 12.20575, 12.82536, 12.94756, 12.22782, 12.36007,
    12.50046, 12.26748, 12.1962, 12.21736, 12.19006, 12.58211, 12.87025,
    12.5106, 12.38481, 12.71254, 12.80705, 12.41378, 14.37295, 15.85056,
    13.81054, 12.82607,
  12.3786, 12.414, 12.24366, 12.46832, 12.36075, 12.22418, 12.24478,
    12.25992, 12.28912, 12.40458, 12.87157, 13.30453, 13.37846, 12.94529,
    12.76674, 12.76902, 12.31042, 12.31284, 12.67011, 13.18279, 13.1995,
    12.56863, 12.33484, 12.82279, 15.8272, 16.43588, 15.97648, 19.38199,
    15.13023, 13.60618,
  12.39539, 12.42015, 12.32804, 12.41543, 12.32507, 12.21749, 12.20549,
    12.26132, 12.35338, 12.41944, 12.48408, 12.85994, 13.22917, 13.50596,
    13.52695, 12.82613, 12.63385, 12.98238, 13.05333, 13.10892, 13.37312,
    14.08991, 14.90241, 14.26384, 18.80875, 22.33643, 18.12399, 19.30304,
    15.02669, 14.09754,
  12.2994, 12.29726, 12.45109, 12.54624, 12.70699, 13.0767, 13.09542,
    12.84558, 12.80704, 12.99218, 13.09229, 13.40667, 13.26483, 13.04212,
    13.76483, 14.35799, 13.90877, 13.0281, 12.84527, 12.69724, 14.64389,
    16.20671, 15.41432, 19.25285, 21.63946, 19.91997, 21.46614, 18.71777,
    14.8989, 13.41655,
  12.62925, 12.37167, 12.56866, 12.82264, 13.13078, 13.37672, 13.27951,
    12.98989, 13.39053, 13.99393, 14.06698, 13.7597, 13.2898, 13.37595,
    14.09284, 14.53941, 13.34722, 12.34077, 12.50982, 16.44849, 18.55964,
    14.83815, 14.59108, 17.24732, 19.01561, 18.35335, 18.37984, 18.4458,
    18.38976, 14.46491,
  12.5637, 12.44814, 13.04008, 14.0273, 14.23929, 13.78611, 13.56346,
    13.27671, 13.12856, 13.30784, 13.15729, 14.26955, 15.89835, 16.16721,
    15.30167, 19.83875, 25.37686, 19.57059, 15.19662, 18.14002, 17.28368,
    13.59645, 14.26394, 14.973, 17.3041, 17.26593, 18.22193, 29.05087,
    27.77213, 14.29531,
  12.4823, 12.70312, 13.5489, 14.68829, 15.1154, 14.49927, 14.39228,
    15.57575, 15.67205, 15.5416, 16.2191, 16.39625, 15.82263, 15.44225,
    19.41303, 27.06, 26.46761, 18.75308, 16.09963, 16.17162, 14.74914,
    13.79555, 14.26025, 16.17064, 17.77572, 15.29116, 23.41937, 40.76498,
    31.13127, 12.85724,
  12.6111, 12.92905, 13.87256, 14.86374, 14.76274, 16.1593, 18.03569,
    16.63528, 15.47024, 15.73451, 16.0022, 15.15621, 13.85386, 13.6604,
    16.76473, 19.88682, 18.15404, 16.07271, 14.91519, 14.70585, 14.25263,
    13.92866, 14.90669, 17.08478, 17.15272, 14.596, 28.97232, 39.06818,
    20.51988, 12.99205,
  13.77641, 13.83317, 14.84166, 15.10388, 15.34971, 18.01534, 17.86132,
    15.46036, 15.43831, 15.73249, 15.08045, 13.99626, 13.3026, 16.38119,
    18.75408, 16.09094, 15.95846, 17.58243, 17.55856, 15.69027, 13.88223,
    14.86571, 18.54053, 19.75724, 16.58618, 16.21187, 24.68985, 25.55471,
    14.7703, 13.21411,
  15.68472, 16.60475, 18.24374, 19.89067, 20.35106, 18.23956, 14.98545,
    14.55164, 14.44464, 13.77176, 14.35271, 17.51154, 19.25239, 19.67539,
    18.90294, 18.37066, 18.92501, 19.82866, 19.44995, 18.07244, 17.54066,
    18.6678, 20.52308, 19.11008, 22.58198, 31.78554, 27.08602, 16.696,
    13.94575, 12.46814,
  22.0402, 25.24599, 24.19415, 20.82692, 20.57887, 20.06524, 17.09928,
    18.32531, 19.12931, 24.28078, 28.23181, 20.15886, 18.12129, 17.66267,
    16.70564, 17.70592, 19.2505, 19.5667, 18.6761, 18.41991, 20.90635,
    21.2232, 18.53708, 16.1002, 20.78105, 26.72893, 20.97804, 13.65709,
    12.80198, 12.17411,
  35.37694, 27.65209, 26.64734, 27.26448, 26.14594, 22.52599, 26.11715,
    25.38538, 20.70534, 25.96248, 27.08811, 16.13591, 16.71766, 18.01629,
    17.1691, 17.60005, 17.26494, 17.39418, 17.16189, 17.779, 21.04768,
    20.31832, 15.77336, 18.70796, 21.76771, 16.44512, 12.99477, 12.94901,
    12.9326, 12.40841,
  49.79226, 39.00592, 42.55935, 49.87831, 51.3404, 47.51443, 37.64668,
    23.09647, 22.50048, 22.71093, 20.16783, 13.89362, 18.59155, 21.80074,
    18.60126, 17.74462, 17.82271, 17.19917, 16.70316, 19.47766, 21.78666,
    18.41123, 15.35328, 21.25278, 24.01217, 14.97772, 12.80916, 13.20019,
    13.51673, 12.78048,
  51.65776, 66.4408, 65.93357, 69.33544, 65.66123, 56.02671, 40.83654,
    36.08981, 29.44522, 25.72301, 31.02894, 30.88946, 34.98657, 35.30449,
    30.87657, 24.18983, 18.31208, 19.7852, 21.23234, 22.83503, 20.78377,
    19.68328, 22.42557, 19.91835, 16.80838, 13.49892, 12.91258, 12.85526,
    13.31945, 12.81449,
  33.87033, 40.69756, 41.78519, 44.56044, 40.77842, 39.46972, 49.19559,
    49.41249, 39.49163, 40.18959, 42.55314, 33.91124, 26.72035, 31.4356,
    34.20125, 22.71664, 21.64159, 21.78546, 23.50266, 25.45655, 23.87523,
    21.73867, 19.67152, 15.80078, 12.97262, 13.4045, 12.98674, 12.69539,
    12.7478, 12.48642,
  22.74277, 23.2515, 25.10139, 25.33248, 23.50516, 27.05582, 34.61721,
    31.96223, 29.69069, 31.79147, 30.84942, 23.9515, 19.34191, 23.97797,
    24.22084, 21.20467, 23.28252, 21.56022, 21.51166, 22.66216, 19.90642,
    17.38094, 14.33603, 13.73841, 13.66233, 13.38296, 13.0263, 12.78955,
    12.62686, 12.35345,
  21.68277, 21.57315, 21.11625, 20.0099, 19.68379, 20.89277, 22.07007,
    21.67702, 22.09412, 22.91689, 20.12292, 20.13252, 23.22786, 21.80666,
    21.41953, 21.84351, 22.20883, 19.96032, 20.41097, 20.44243, 15.07066,
    14.63915, 14.19664, 13.90187, 13.56701, 13.44058, 12.99114, 12.57597,
    12.53918, 12.35328,
  19.51166, 19.03052, 17.90654, 17.82591, 18.27115, 19.3456, 20.23723,
    20.75789, 20.74505, 19.16768, 18.69175, 22.63583, 24.69601, 23.60932,
    25.89532, 24.53501, 20.70777, 17.69872, 19.88395, 19.41779, 14.35863,
    14.40087, 14.26483, 13.98573, 13.20765, 13.17571, 12.9453, 12.38394,
    12.3573, 12.25882,
  19.28596, 18.95952, 17.38062, 16.95416, 17.49285, 18.10775, 18.65905,
    18.82308, 18.09301, 17.19534, 20.05599, 22.5002, 20.40869, 21.45358,
    23.09088, 21.86833, 20.50467, 19.55377, 21.43215, 20.40472, 16.63277,
    15.29043, 14.36402, 14.01428, 13.03505, 12.82217, 12.76076, 12.37613,
    12.29115, 12.21521,
  19.57613, 19.33252, 17.84456, 16.64033, 16.97847, 17.1039, 17.16524,
    17.087, 16.71249, 18.80185, 21.59012, 19.88437, 18.14012, 18.63888,
    18.60748, 17.96247, 18.78061, 20.23508, 21.02605, 21.16305, 19.70029,
    17.09332, 14.47166, 14.04394, 13.32413, 12.8198, 12.66353, 12.40525,
    12.28911, 12.21687,
  19.01054, 19.1121, 17.82851, 16.63084, 16.5775, 16.61523, 16.50908,
    16.43813, 17.26918, 20.37312, 20.76199, 17.57711, 17.96518, 17.96451,
    17.07388, 16.30875, 16.52299, 17.23276, 17.84487, 18.35154, 18.84687,
    18.20191, 15.80471, 14.61911, 13.80194, 13.12329, 12.64731, 12.39963,
    12.29014, 12.21475,
  19.67532, 18.91484, 17.70657, 16.93497, 16.73875, 16.26709, 16.37783,
    16.71729, 18.56928, 20.78138, 18.99751, 16.37058, 17.06368, 16.91413,
    16.19156, 15.77008, 15.47649, 15.33445, 15.80257, 15.92022, 17.04106,
    17.3898, 16.02011, 16.35029, 15.13647, 13.4692, 12.70952, 12.47607,
    12.29059, 12.21305,
  19.87168, 19.08314, 17.57244, 16.75381, 17.18452, 17.4966, 17.80602,
    17.72713, 19.25186, 19.88163, 17.22733, 15.87163, 16.08176, 15.91794,
    15.39263, 15.63144, 15.63734, 14.8933, 14.69769, 14.66712, 15.91406,
    15.92504, 14.39526, 16.04213, 16.23808, 14.16051, 12.90594, 12.90777,
    12.59695, 12.25046,
  19.64408, 19.0341, 18.08682, 17.87702, 18.48495, 18.93444, 20.11096,
    20.84426, 21.54161, 19.34957, 16.22641, 16.09247, 16.25752, 16.37784,
    16.02061, 16.10484, 16.29054, 15.38209, 14.45788, 14.582, 15.03331,
    14.6304, 13.8885, 14.39054, 15.3704, 15.49796, 14.27687, 13.35605,
    13.07028, 12.42928,
  19.65303, 19.57879, 18.23416, 18.22044, 19.4027, 20.13782, 20.42429,
    20.73735, 21.76123, 19.483, 15.97737, 16.24045, 16.50903, 16.69967,
    16.62617, 16.64319, 16.28237, 15.75467, 15.02972, 14.63513, 14.57249,
    14.3798, 14.29618, 13.88739, 13.899, 15.35355, 15.63252, 14.34345,
    14.02186, 12.95492,
  19.95473, 20.90946, 20.41735, 19.9862, 20.07621, 20.07291, 20.62378,
    21.55304, 20.57753, 18.38351, 16.27022, 16.57783, 17.01681, 16.74142,
    16.18421, 16.14043, 15.75193, 15.60485, 15.48098, 14.8687, 14.76262,
    14.7716, 14.1132, 13.53032, 13.52034, 14.37554, 15.92496, 15.16968,
    14.07865, 12.99247,
  21.08292, 22.28592, 21.52333, 20.70822, 19.98227, 19.19785, 20.96129,
    21.81011, 18.97358, 16.77221, 16.64729, 17.13991, 17.26008, 16.61787,
    15.85686, 15.48766, 15.26802, 15.40809, 15.35437, 14.70928, 14.7222,
    15.53633, 15.5463, 14.95892, 15.05112, 15.4139, 17.43045, 17.12006,
    13.98303, 12.38655,
  22.12805, 22.85253, 20.76956, 20.4165, 20.53582, 19.85495, 20.86976,
    20.09928, 16.8514, 16.12724, 16.59628, 16.97115, 16.79543, 16.31025,
    16.17511, 15.75072, 15.12066, 15.03242, 15.48973, 15.88417, 16.16997,
    16.33024, 16.04812, 15.66177, 15.92718, 16.16656, 16.95101, 18.76276,
    16.75972, 12.99891,
  21.04889, 20.22748, 20.22313, 21.84583, 22.25203, 22.0234, 21.28677,
    18.32467, 16.09031, 16.26877, 15.94481, 15.52642, 15.36142, 15.40378,
    15.89258, 16.0166, 15.83677, 16.15952, 16.253, 16.06662, 16.09851,
    15.70081, 14.83804, 14.44834, 14.85108, 15.42021, 15.58861, 15.98787,
    16.49577, 13.8306,
  20.36948, 20.0366, 20.4214, 21.04116, 21.08075, 22.1856, 21.83319,
    18.17289, 15.93964, 16.29366, 16.26672, 16.33478, 16.52664, 16.74675,
    16.95828, 17.05038, 16.48605, 15.73913, 15.44709, 14.79888, 14.26267,
    14.16771, 13.89471, 13.7357, 13.91234, 14.54067, 14.76681, 14.07722,
    13.66404, 12.70271,
  13.19964, 13.22412, 13.2556, 13.26752, 13.26369, 13.25896, 13.2469,
    13.26156, 13.28517, 13.27378, 13.9042, 14.05182, 13.28361, 13.43009,
    13.59267, 13.36651, 13.3012, 13.31728, 13.28429, 13.68462, 13.98654,
    13.60664, 13.48851, 13.81807, 13.87965, 13.45221, 15.41354, 17.10814,
    15.01307, 14.00086,
  13.45735, 13.5065, 13.32479, 13.55765, 13.45314, 13.30654, 13.32721,
    13.34116, 13.36556, 13.4852, 14.01845, 14.45343, 14.45616, 14.05934,
    13.8604, 13.88326, 13.42063, 13.40549, 13.77191, 14.36395, 14.4087,
    13.70776, 13.40353, 13.88519, 16.81927, 17.67366, 17.21429, 21.17933,
    16.48479, 14.82369,
  13.49076, 13.51547, 13.42147, 13.52915, 13.42982, 13.29821, 13.2717,
    13.34476, 13.44343, 13.52603, 13.60304, 14.00419, 14.43189, 14.68309,
    14.683, 13.9504, 13.7172, 14.08543, 14.21411, 14.32118, 14.54555,
    15.18985, 15.94654, 15.25386, 19.76515, 24.05527, 19.61132, 21.18567,
    16.37026, 15.38384,
  13.37966, 13.36177, 13.51681, 13.61494, 13.78548, 14.19773, 14.19772,
    13.93352, 13.90574, 14.07983, 14.21478, 14.60415, 14.46471, 14.18465,
    14.94518, 15.56415, 15.1802, 14.23946, 13.99719, 13.75813, 15.72796,
    17.44753, 16.52692, 20.20868, 23.00855, 21.5728, 23.42457, 20.63397,
    16.33534, 14.68561,
  13.72026, 13.45369, 13.62835, 13.86939, 14.2485, 14.57883, 14.4537,
    14.10737, 14.52312, 15.23902, 15.39621, 15.05781, 14.43469, 14.44022,
    15.29804, 15.8757, 14.65692, 13.44322, 13.51488, 17.32225, 19.83118,
    16.07471, 15.63562, 18.46552, 20.4447, 19.81104, 20.2152, 20.25105,
    20.02868, 15.78467,
  13.67501, 13.52269, 14.10154, 15.10201, 15.42626, 15.01716, 14.72037,
    14.41636, 14.31038, 14.58246, 14.39343, 15.40408, 17.121, 17.42158,
    16.5848, 20.93501, 26.62979, 20.77212, 16.23956, 19.38105, 18.72267,
    14.62956, 15.33938, 16.16796, 18.68872, 18.8979, 19.40464, 31.03154,
    30.67648, 15.71425,
  13.56085, 13.77026, 14.63991, 15.81415, 16.30897, 15.73725, 15.64095,
    17.02021, 17.08965, 16.81248, 17.3849, 17.63232, 17.23982, 16.80784,
    20.75193, 29.18251, 28.91005, 20.31764, 17.37139, 17.51592, 15.88774,
    14.81622, 15.40136, 17.51878, 19.37723, 16.82248, 24.13448, 43.19628,
    35.24752, 14.22184,
  13.67432, 14.01153, 14.96589, 15.98702, 15.91614, 17.37752, 19.61232,
    18.39871, 17.02202, 17.16525, 17.45062, 16.55445, 15.06122, 14.77583,
    18.24204, 22.09646, 19.97883, 17.36084, 16.09701, 15.88348, 15.35994,
    15.01225, 16.07164, 18.55532, 18.68966, 15.87855, 30.03296, 42.19329,
    23.36342, 14.25202,
  14.83914, 14.92329, 15.93387, 16.20911, 16.47083, 19.58555, 19.77751,
    16.94528, 16.73065, 17.12911, 16.43366, 15.12969, 14.28191, 17.48448,
    20.21603, 17.41519, 17.22706, 18.98468, 18.86539, 16.96638, 14.99993,
    15.96482, 19.84542, 21.36659, 17.88992, 17.38013, 26.56298, 28.37746,
    16.16184, 14.44279,
  16.98022, 17.66557, 19.54155, 21.68459, 22.00212, 19.9391, 16.36906,
    15.79278, 15.77122, 15.12901, 15.45136, 18.51361, 20.34308, 21.14514,
    20.54094, 19.69869, 20.27169, 21.33228, 21.01101, 19.40792, 18.77336,
    19.93673, 22.06595, 20.6223, 22.98407, 32.23593, 29.04563, 18.50205,
    15.26135, 13.6395,
  22.32349, 26.29877, 26.14991, 22.483, 22.17013, 21.71514, 18.50116,
    19.72189, 20.60853, 24.66041, 28.88721, 21.7455, 19.57783, 19.07577,
    18.03601, 19.09073, 20.80389, 21.11509, 20.201, 19.78899, 22.42788,
    22.90364, 20.09768, 17.1955, 21.66643, 28.37753, 23.17935, 14.99356,
    13.97372, 13.2895,
  37.13455, 29.45513, 27.4315, 26.9624, 26.20812, 22.41343, 26.82828,
    27.30516, 22.12967, 26.83327, 28.49125, 17.54151, 17.84456, 19.12302,
    18.44547, 19.05859, 18.72751, 18.85032, 18.5113, 19.12714, 22.72915,
    22.10026, 17.05508, 19.58224, 23.12089, 18.15669, 14.36451, 14.0982,
    14.10015, 13.52754,
  50.6793, 37.12074, 40.2111, 47.2697, 50.59524, 48.85076, 41.14542,
    24.88817, 24.48687, 24.31494, 21.35365, 14.9935, 19.84869, 23.08781,
    19.97958, 19.05019, 19.24298, 18.58069, 18.00243, 21.07223, 23.82293,
    20.01785, 16.49232, 22.54787, 26.22074, 16.5806, 13.95351, 14.34499,
    14.72686, 13.97204,
  53.13555, 58.43523, 58.12004, 63.65707, 65.12361, 60.78323, 45.03991,
    37.80801, 31.32266, 26.351, 31.28185, 31.36688, 36.4684, 36.77868,
    32.45799, 25.62468, 19.76803, 21.38556, 23.13389, 25.23738, 22.94326,
    20.77645, 23.80251, 22.07487, 18.94092, 14.84162, 14.05652, 14.01863,
    14.53064, 14.00956,
  35.33111, 38.65935, 41.95438, 51.15124, 53.56347, 46.99089, 49.49801,
    49.8749, 39.22335, 39.79454, 42.95214, 35.51792, 28.9928, 34.01626,
    36.92418, 24.77123, 23.46244, 23.80612, 25.86791, 27.76966, 25.32186,
    23.32264, 21.83355, 17.88207, 14.24064, 14.60786, 14.15179, 13.83118,
    13.89716, 13.64124,
  23.70008, 25.76346, 30.8829, 35.03206, 32.88848, 30.65365, 35.30509,
    32.38665, 30.00402, 32.93748, 32.54112, 25.6599, 20.58398, 26.08604,
    26.68931, 23.20049, 25.69511, 23.84002, 23.50635, 24.71496, 21.72828,
    19.39173, 16.1484, 15.19721, 14.87823, 14.57345, 14.18886, 13.92913,
    13.74958, 13.47157,
  22.36574, 23.55548, 24.24674, 22.7949, 20.76898, 21.21169, 22.66224,
    22.00061, 22.65248, 23.96662, 21.09347, 20.92567, 24.32439, 23.26468,
    23.31824, 23.96784, 24.68, 22.13273, 22.23633, 22.73741, 17.00674,
    16.35284, 15.60979, 15.19167, 14.77345, 14.6291, 14.15941, 13.72656,
    13.66051, 13.46581,
  19.89068, 19.81426, 18.34684, 17.51099, 17.64069, 18.93417, 19.94557,
    20.65065, 20.8807, 19.253, 18.68544, 23.18682, 25.94462, 24.88146,
    28.37683, 27.32949, 23.08913, 19.55245, 21.95856, 21.92178, 16.12631,
    15.94969, 15.56789, 15.25054, 14.41782, 14.36926, 14.12916, 13.51225,
    13.47417, 13.37656,
  19.42707, 18.95188, 16.94707, 16.31901, 16.85476, 17.5098, 18.16323,
    18.47978, 17.80424, 16.6519, 19.80207, 23.06023, 21.21918, 22.76927,
    25.65656, 24.62248, 22.92126, 21.51575, 23.68212, 22.64515, 18.20881,
    16.64711, 15.66052, 15.32657, 14.25769, 14.00373, 13.94841, 13.50827,
    13.40339, 13.32052,
  19.58599, 18.96327, 17.16023, 15.81376, 16.19541, 16.39849, 16.60186,
    16.58952, 16.02637, 18.06889, 21.47581, 20.23561, 18.59382, 19.81628,
    20.50946, 20.06871, 21.07482, 22.58188, 23.2043, 23.26517, 21.49859,
    18.66836, 15.83341, 15.37183, 14.57195, 14.01182, 13.82665, 13.54121,
    13.40709, 13.32888,
  18.75838, 18.54112, 17.11486, 15.79731, 15.82808, 15.98404, 15.91074,
    15.68973, 16.38012, 19.87829, 20.90144, 17.76048, 18.61831, 19.21313,
    18.72379, 18.14101, 18.5298, 19.21946, 19.58582, 20.20338, 20.77796,
    20.03108, 17.23368, 15.93218, 15.05343, 14.34494, 13.82446, 13.54471,
    13.40324, 13.32501,
  19.27207, 18.25235, 17.00283, 16.17776, 16.06272, 15.5995, 15.60357,
    15.81697, 17.83524, 20.59275, 19.0979, 16.56377, 17.89472, 18.29423,
    17.86817, 17.50609, 17.20427, 16.84988, 17.33457, 17.54493, 18.75642,
    19.30754, 17.50575, 17.73736, 16.5013, 14.75687, 13.86935, 13.60928,
    13.4, 13.32366,
  19.39339, 18.40705, 16.91226, 16.08558, 16.56971, 16.75301, 16.95433,
    16.87959, 18.80443, 19.94129, 17.26177, 16.19233, 17.02109, 17.32367,
    17.00634, 17.29521, 17.21765, 16.31881, 16.14666, 16.10513, 17.56112,
    17.76385, 15.74558, 17.62277, 17.89095, 15.54474, 14.04822, 14.04625,
    13.68362, 13.34784,
  19.1802, 18.44448, 17.47804, 17.13448, 17.69995, 18.13951, 19.48966,
    20.55806, 21.58991, 19.46823, 16.23024, 16.56552, 17.25448, 17.77194,
    17.57365, 17.68041, 17.87413, 16.91516, 15.86774, 15.92701, 16.59026,
    16.20144, 15.16747, 15.85763, 17.01873, 16.97509, 15.54415, 14.54043,
    14.159, 13.52479,
  19.23929, 19.16373, 17.63964, 17.36878, 18.55827, 19.48954, 20.14859,
    20.93315, 22.22895, 19.81547, 16.08335, 16.76986, 17.53609, 18.09326,
    18.17977, 18.30606, 17.96505, 17.36153, 16.42334, 15.9745, 15.92663,
    15.64154, 15.58802, 15.22745, 15.22583, 16.74737, 16.99391, 15.55385,
    15.17124, 14.119,
  19.56321, 20.42349, 19.68876, 19.16657, 19.40167, 19.76578, 20.62025,
    21.89451, 21.00325, 18.73105, 16.36325, 16.94341, 17.88817, 18.0866,
    17.76299, 17.8887, 17.45024, 17.1342, 16.86817, 16.14208, 16.00989,
    16.05225, 15.41583, 14.79107, 14.70478, 15.59635, 17.19209, 16.4669,
    15.37063, 14.23358,
  20.68951, 21.55199, 20.83911, 20.05574, 19.48698, 18.98507, 21.25691,
    22.5507, 19.32802, 16.85044, 16.64964, 17.42001, 18.08249, 17.92672,
    17.38598, 17.0773, 16.81572, 16.87546, 16.76577, 16.0216, 15.99607,
    16.86027, 16.88825, 16.19177, 16.21826, 16.58048, 18.68905, 18.46952,
    15.24876, 13.56872,
  21.81162, 22.37158, 20.10159, 19.91324, 20.23957, 19.88812, 21.34765,
    20.77798, 16.98475, 15.96028, 16.54732, 17.32059, 17.62684, 17.55416,
    17.60252, 17.21931, 16.55834, 16.45654, 16.8393, 17.23246, 17.61495,
    17.81215, 17.51762, 17.03238, 17.16024, 17.45843, 18.38381, 20.27815,
    18.18034, 14.17713,
  20.72019, 19.70283, 19.74443, 21.84621, 22.49286, 22.54766, 22.11944,
    18.80468, 15.97439, 16.06146, 15.94297, 15.94823, 16.18754, 16.54931,
    17.29785, 17.48851, 17.25487, 17.60668, 17.66945, 17.57719, 17.69851,
    17.18061, 16.19462, 15.73469, 16.10266, 16.69993, 16.91806, 17.52207,
    18.01982, 15.11136,
  20.11811, 19.73272, 20.51499, 21.4909, 21.6842, 23.06708, 22.7712,
    18.50545, 15.80599, 16.23387, 16.35175, 16.6766, 17.20207, 17.7501,
    18.21839, 18.4571, 17.94075, 17.28763, 16.93968, 16.19366, 15.60673,
    15.45918, 15.11954, 14.92729, 15.11586, 15.75599, 16.04938, 15.33216,
    14.9426, 13.93466,
  19.0074, 19.06248, 19.07035, 19.08564, 19.0818, 19.07447, 19.06305,
    19.10066, 19.131, 19.15284, 19.96434, 20.20123, 19.16795, 19.33566,
    19.55218, 19.2466, 19.13734, 19.17472, 19.17364, 19.72535, 20.15556,
    19.63191, 19.50723, 19.86621, 19.9301, 19.50656, 21.83376, 24.36022,
    21.59483, 20.25629,
  19.31097, 19.43326, 19.14355, 19.44257, 19.30878, 19.12451, 19.14251,
    19.18711, 19.24004, 19.41422, 20.07987, 20.67117, 20.73346, 20.20639,
    19.86906, 19.91683, 19.30304, 19.30836, 19.8545, 20.68415, 20.66442,
    19.70252, 19.32149, 19.97418, 23.45506, 25.36414, 24.44976, 30.09792,
    23.68363, 21.44312,
  19.37317, 19.40797, 19.27255, 19.40922, 19.30257, 19.14001, 19.09751,
    19.20724, 19.35036, 19.46976, 19.62251, 20.15602, 20.65587, 20.95725,
    20.98527, 20.01304, 19.73722, 20.28067, 20.43683, 20.58308, 20.90958,
    21.88206, 22.76576, 22.0809, 26.83455, 32.77903, 27.94404, 30.17998,
    23.5614, 22.27923,
  19.25002, 19.23931, 19.41583, 19.5562, 19.79877, 20.30641, 20.33118,
    20.01771, 19.98056, 20.19318, 20.37957, 20.88736, 20.73875, 20.30745,
    21.39158, 22.32002, 21.83682, 20.50077, 20.09477, 19.89747, 22.44192,
    24.84445, 23.56106, 28.02736, 31.60761, 29.57225, 33.23455, 29.07079,
    23.4094, 21.21328,
  19.74072, 19.35095, 19.59446, 19.92741, 20.39055, 20.77917, 20.66598,
    20.26065, 20.78484, 21.82129, 22.10022, 21.47039, 20.58274, 20.85292,
    22.05475, 22.61618, 21.109, 19.39517, 19.5968, 24.45245, 28.06939,
    22.88041, 22.40345, 25.64547, 28.15692, 27.62588, 28.32605, 29.1817,
    28.96599, 22.64849,
  19.66028, 19.46125, 20.23772, 21.55203, 21.99903, 21.44179, 20.97664,
    20.63393, 20.49475, 20.86094, 20.67402, 21.8747, 24.19532, 24.60015,
    23.94575, 28.91841, 36.29088, 29.35953, 23.39179, 27.01614, 26.17383,
    20.97708, 21.85732, 23.09964, 26.09199, 26.55535, 26.61126, 41.04791,
    42.25331, 22.51678,
  19.50239, 19.79264, 20.88626, 22.362, 23.04838, 22.38215, 22.12345,
    23.97169, 24.1179, 23.79632, 24.51876, 24.83347, 24.27071, 23.89524,
    28.6281, 38.52362, 38.22554, 28.20207, 24.58289, 24.6721, 22.55788,
    21.13946, 21.88186, 24.58414, 26.90607, 24.27431, 31.53871, 52.82912,
    45.91833, 20.75945,
  19.627, 20.10452, 21.29732, 22.57059, 22.48452, 24.20514, 27.16421,
    25.80581, 23.95529, 24.23025, 24.51344, 23.42843, 21.51534, 21.41159,
    25.68738, 30.21879, 27.42097, 24.63867, 22.86525, 22.54956, 21.81222,
    21.32156, 22.72172, 25.86951, 26.06744, 23.31608, 38.37149, 53.05576,
    31.5819, 20.60394,
  21.19707, 21.35642, 22.43745, 22.67646, 23.15229, 27.49832, 27.90594,
    23.90652, 23.78569, 24.2877, 23.36102, 21.61567, 20.64579, 24.68483,
    28.67798, 25.13854, 24.30829, 26.51131, 26.41966, 24.04691, 21.35159,
    22.64572, 27.52082, 29.6145, 25.06084, 24.84985, 35.15022, 37.97521,
    23.40933, 20.68425,
  23.56555, 24.14776, 26.73475, 30.3135, 30.53738, 28.0188, 23.23097,
    22.36953, 22.35748, 21.68771, 21.9661, 25.77143, 28.12835, 29.22775,
    28.35749, 27.3819, 28.33511, 29.5203, 28.90339, 26.83553, 26.16003,
    27.40032, 29.93114, 28.57433, 31.58313, 43.10854, 39.55176, 25.91013,
    21.6057, 19.62719,
  31.70112, 37.41734, 37.86435, 30.39651, 30.40618, 30.3208, 26.90509,
    27.88068, 29.16736, 32.71808, 38.03028, 29.8526, 27.35896, 26.73347,
    25.55119, 26.93111, 29.27206, 29.66953, 28.25242, 27.11839, 30.32921,
    30.83162, 27.39646, 24.13317, 29.53838, 37.52691, 31.36879, 21.20107,
    20.07528, 19.13276,
  48.53906, 40.09987, 36.60087, 33.90395, 34.49944, 29.79296, 34.58978,
    34.908, 29.96946, 35.02332, 36.49243, 23.98192, 24.92365, 26.68682,
    25.91515, 26.90858, 26.6477, 26.73711, 26.04932, 26.50729, 30.80588,
    29.89449, 23.71113, 26.57501, 31.48338, 25.73627, 20.76489, 20.20507,
    20.18025, 19.44672,
  61.41715, 47.96243, 50.73546, 57.35763, 59.02878, 56.29959, 50.47198,
    43.55322, 49.47869, 36.42939, 27.54478, 22.63341, 28.5732, 30.70264,
    28.44717, 26.6762, 27.01546, 26.07815, 25.06078, 28.75805, 32.22147,
    27.16548, 23.05274, 29.89656, 35.00088, 23.36213, 20.04863, 20.51837,
    20.92138, 20.00838,
  69.8268, 60.43312, 62.31311, 67.96791, 71.15622, 71.60945, 63.12409,
    61.27783, 51.53181, 36.06461, 40.15281, 42.4751, 48.30615, 49.46622,
    43.26812, 33.43097, 27.78152, 29.78296, 32.05458, 34.89291, 31.76212,
    27.69735, 32.13217, 30.15442, 26.19741, 21.234, 20.18001, 20.13026,
    20.69705, 20.09543,
  53.06149, 63.84921, 72.33765, 79.62495, 80.39795, 70.70007, 67.98586,
    69.27313, 48.97008, 49.55314, 57.27216, 49.18126, 40.31614, 42.62371,
    47.89433, 33.71286, 32.64368, 33.23564, 35.94133, 38.0147, 33.51347,
    30.99334, 29.89335, 25.2365, 20.61757, 20.96505, 20.33887, 19.93143,
    19.93851, 19.61733,
  39.37984, 49.25608, 56.43069, 55.88683, 49.34472, 49.56389, 53.86641,
    41.54063, 43.15018, 49.9242, 41.85892, 37.19346, 29.41565, 34.00387,
    35.47298, 32.25685, 35.7478, 33.3383, 32.18431, 33.55523, 29.23097,
    26.48025, 23.11501, 21.79705, 21.27014, 20.90469, 20.38449, 20.04044,
    19.75578, 19.39202,
  31.1486, 32.54861, 33.08035, 29.47924, 26.80168, 30.93163, 33.49361,
    29.12339, 34.00486, 36.12247, 27.06945, 27.91678, 31.83183, 30.73659,
    31.3416, 32.68316, 34.28234, 30.98261, 30.3018, 31.81639, 24.11932,
    23.00751, 22.07237, 21.72289, 21.15216, 20.89436, 20.33183, 19.76042,
    19.61217, 19.38501,
  24.67482, 24.72848, 22.6078, 21.41025, 22.00421, 24.03495, 25.35396,
    26.46207, 26.59303, 24.12202, 23.1814, 28.69497, 32.86319, 31.8421,
    37.85815, 36.94328, 31.81027, 27.21815, 30.20535, 30.6986, 22.73595,
    22.6341, 22.13542, 21.79336, 20.65469, 20.56892, 20.31576, 19.48208,
    19.3922, 19.26287,
  23.64263, 22.98227, 20.0639, 19.21765, 20.03094, 20.94379, 21.96438,
    22.28893, 21.19267, 19.51456, 23.38294, 27.93103, 26.10379, 29.0035,
    34.3875, 33.32718, 31.41083, 29.4177, 32.44363, 31.1137, 25.25699,
    23.53976, 22.32311, 21.89652, 20.46633, 20.14562, 20.06375, 19.44804,
    19.32171, 19.2134,
  23.44526, 22.31891, 19.77625, 18.05542, 18.6292, 18.95944, 19.22254,
    19.18643, 18.3827, 20.82231, 25.35444, 23.9467, 22.3368, 25.13721,
    27.27153, 27.54801, 29.16466, 31.26075, 31.94211, 31.90948, 29.38427,
    26.07162, 22.64396, 22.00252, 20.90503, 20.16951, 19.90541, 19.51482,
    19.31075, 19.20783,
  21.99939, 21.42698, 19.38422, 17.72807, 17.79254, 17.9987, 17.92691,
    17.62377, 18.43176, 22.84241, 24.39425, 20.41895, 22.22074, 24.11862,
    24.56157, 24.77864, 25.92164, 27.31331, 27.68984, 28.3681, 29.06451,
    28.48383, 24.5252, 22.76948, 21.44331, 20.57287, 19.89628, 19.53895,
    19.32329, 19.21602,
  22.64113, 20.67419, 19.05874, 18.04243, 17.96059, 17.31652, 17.3086,
    17.51544, 20.10543, 23.67059, 21.82433, 18.76002, 21.28516, 22.82132,
    23.40243, 23.90748, 24.21896, 24.14879, 24.8091, 25.08138, 26.67404,
    27.88264, 24.88992, 25.08306, 23.36646, 21.20655, 20.01292, 19.64696,
    19.32492, 19.22456,
  22.63407, 20.68536, 18.83842, 17.82552, 18.5268, 18.7236, 18.8511,
    18.66848, 21.10933, 22.74037, 19.3654, 18.26532, 20.06393, 21.52021,
    22.35663, 23.75712, 24.34561, 23.43808, 23.21206, 23.11936, 24.88776,
    25.70121, 22.74693, 25.04295, 25.29901, 22.29305, 20.19966, 20.18566,
    19.68905, 19.25683,
  22.26176, 20.63794, 19.54516, 19.16498, 19.90716, 20.28384, 22.0197,
    23.70729, 24.99542, 22.09136, 18.02618, 18.69132, 20.30876, 22.1117,
    23.16247, 24.34894, 25.20794, 24.1499, 22.77859, 22.94939, 24.05151,
    23.57129, 21.84793, 22.92698, 24.28368, 24.03361, 22.19038, 20.79326,
    20.24697, 19.4975,
  21.99954, 21.87799, 19.84055, 19.20645, 20.77489, 22.2929, 23.26335,
    24.39579, 25.65293, 22.50488, 17.8415, 19.03274, 20.73165, 22.62662,
    23.96437, 25.21259, 25.31355, 24.6729, 23.44379, 22.92002, 23.0867,
    22.57086, 22.41967, 22.15823, 21.87782, 23.6176, 23.89722, 21.97958,
    21.45271, 20.32878,
  22.51161, 23.79634, 22.6272, 21.69697, 22.03478, 22.84931, 24.19255,
    25.8509, 24.18841, 21.33726, 18.31577, 19.39039, 21.27657, 22.71392,
    23.47156, 24.65798, 24.66784, 24.35059, 23.92948, 22.89042, 22.80857,
    22.99172, 22.27005, 21.32819, 20.97061, 22.05948, 23.85511, 23.1153,
    21.7589, 20.51134,
  23.93648, 25.15521, 24.16891, 22.63041, 22.1203, 21.97634, 25.47629,
    27.18885, 22.38435, 19.19357, 18.89512, 20.10087, 21.61043, 22.48017,
    23.03, 23.69486, 23.84787, 23.97587, 23.7695, 22.71578, 22.83321,
    23.97015, 23.89798, 22.74838, 22.64119, 23.15149, 25.48363, 25.50773,
    21.66921, 19.60563,
  26.14611, 28.01061, 22.81905, 22.07006, 22.90728, 23.01565, 25.32899,
    24.81942, 19.60307, 18.23598, 19.01709, 20.17761, 21.09914, 21.90635,
    23.30318, 23.91184, 23.47961, 23.4357, 23.76777, 23.97598, 24.6698,
    25.28104, 24.77222, 23.93031, 23.82862, 24.29595, 25.4653, 27.71793,
    25.32213, 20.35413,
  24.57035, 23.08911, 22.27748, 26.54144, 27.11028, 26.16649, 26.15365,
    22.12164, 18.3068, 18.45309, 18.3624, 18.47895, 19.1905, 20.54331,
    22.73052, 24.09448, 24.2548, 24.81395, 24.86104, 24.47002, 24.78916,
    24.35945, 23.04066, 22.32344, 22.69925, 23.48889, 23.93817, 24.81409,
    25.1195, 21.58634,
  23.31573, 22.30218, 24.4586, 27.63517, 27.19911, 27.66482, 27.30163,
    22.02266, 18.25966, 18.89503, 18.97667, 19.37619, 20.43996, 21.98252,
    23.73715, 25.02408, 24.98443, 24.46959, 23.97838, 22.89218, 22.18324,
    21.94254, 21.50604, 21.22232, 21.53252, 22.36255, 22.83128, 22.07118,
    21.42159, 20.09272,
  16.66882, 16.76019, 16.8028, 16.8613, 16.86471, 16.86592, 16.86176,
    16.91225, 16.97026, 17.25399, 18.88377, 19.3731, 17.1807, 17.5154, 17.86,
    17.18664, 16.95905, 16.99912, 17.17176, 18.11915, 18.68286, 18.21278,
    18.52986, 19.30007, 20.03992, 20.48738, 24.96012, 29.22858, 21.85333,
    18.90047,
  17.41735, 17.6473, 17.07705, 17.63106, 17.35573, 17.02601, 17.10948,
    17.22195, 17.43978, 17.936, 19.01214, 20.0783, 20.40737, 19.29541,
    18.41542, 18.60329, 17.45332, 17.66328, 18.88684, 20.14202, 19.5341,
    18.25032, 18.89898, 22.11504, 29.67895, 33.64703, 30.39311, 37.09604,
    24.47532, 20.5099,
  17.36517, 17.41157, 17.2377, 17.37635, 17.16194, 16.99087, 17.05369,
    17.28122, 17.55877, 17.76585, 18.09031, 19.04583, 19.83184, 20.51708,
    20.65825, 18.82077, 18.7287, 19.7767, 19.84175, 20.30223, 21.95005,
    25.6017, 28.49022, 30.32956, 39.65701, 46.38807, 37.79693, 37.0822,
    24.68259, 21.95615,
  17.2083, 17.26999, 17.60599, 17.95436, 18.42476, 19.34706, 19.45158,
    18.86946, 18.84388, 19.43421, 19.98706, 20.50055, 20.17649, 19.61922,
    21.80276, 23.67282, 22.69481, 20.12223, 19.93694, 21.46159, 27.70725,
    32.52715, 30.7178, 39.02656, 46.59315, 40.88586, 45.4998, 35.12238,
    24.49496, 19.91055,
  18.14087, 17.52482, 18.1356, 18.78106, 19.62028, 20.01022, 19.72566,
    19.38614, 20.73304, 22.34878, 21.92419, 20.81793, 20.15343, 21.03106,
    22.70751, 23.22935, 21.28824, 19.50679, 22.12018, 31.36937, 36.94276,
    28.18279, 28.91004, 33.5158, 35.81644, 34.85297, 34.41486, 37.69435,
    34.83789, 21.86563,
  18.02787, 18.26675, 19.96394, 22.60313, 22.69727, 20.679, 20.43788,
    20.13076, 19.92743, 20.20458, 20.38032, 23.62426, 28.93883, 29.98632,
    33.38919, 40.80762, 46.43428, 38.95366, 31.41282, 35.29108, 31.97852,
    24.3008, 26.51525, 29.44119, 32.72747, 33.37785, 38.01771, 56.76304,
    51.03709, 20.87794,
  18.33081, 19.589, 21.71118, 23.9104, 23.91934, 22.52272, 24.03451,
    28.11505, 28.59332, 28.65614, 30.48022, 30.57193, 28.99359, 30.56758,
    39.53232, 51.50541, 47.96065, 37.57866, 30.51389, 29.89486, 25.95563,
    23.69042, 25.7484, 30.98089, 35.46886, 38.84994, 50.80702, 64.19802,
    52.04013, 18.7434,
  19.04312, 20.68465, 23.18113, 25.03317, 24.27852, 28.02946, 34.95468,
    32.43009, 28.69744, 29.39222, 28.94026, 27.10387, 25.1676, 27.84599,
    33.89703, 38.10115, 34.81297, 31.32581, 25.76105, 25.14204, 23.64715,
    23.21168, 26.98734, 32.99939, 35.04989, 37.58341, 53.73264, 62.41235,
    37.47964, 18.95271,
  22.19251, 22.92469, 24.93863, 25.89435, 28.52463, 34.7993, 32.93208,
    28.46701, 29.02774, 29.14262, 27.23521, 24.95911, 25.60255, 34.76176,
    41.86797, 33.34841, 30.31036, 33.29872, 33.20193, 28.23152, 23.10067,
    27.46375, 37.18013, 40.90584, 32.99403, 38.84211, 54.4669, 47.33813,
    26.02726, 19.10845,
  28.06281, 33.29659, 36.38596, 39.90901, 42.27308, 38.48759, 25.29627,
    25.06557, 24.44485, 24.89091, 28.58009, 38.17116, 42.93218, 41.39542,
    36.43342, 35.18602, 37.04189, 38.1984, 34.91934, 29.86995, 30.17816,
    32.85154, 36.09285, 37.58302, 47.5811, 62.20938, 52.77482, 27.3862,
    20.02869, 17.32766,
  44.61658, 50.4859, 51.66894, 48.13435, 47.45038, 40.79604, 32.55792,
    36.10798, 40.835, 48.47905, 55.94029, 42.16919, 36.10082, 33.57296,
    31.44125, 33.58038, 36.28226, 35.45054, 32.10843, 29.88863, 33.8477,
    34.62711, 30.02553, 28.0907, 36.38763, 42.90015, 31.36242, 18.53001,
    17.9064, 16.6921,
  66.70457, 53.48882, 53.98492, 55.00558, 52.11671, 43.02742, 51.19149,
    52.84848, 48.53288, 50.93744, 47.26915, 32.32761, 33.19672, 34.98043,
    33.57398, 34.50509, 33.09357, 31.5749, 29.79661, 31.07772, 34.41589,
    31.9271, 24.68637, 29.85001, 36.23011, 26.20961, 18.62533, 18.29447,
    18.14272, 17.11656,
  80.5445, 68.62938, 81.99249, 89.57397, 90.69674, 84.63601, 71.42822,
    54.33691, 55.29677, 44.75378, 36.74937, 31.41387, 40.20142, 45.97524,
    40.82156, 35.17299, 33.67466, 30.80494, 29.20768, 36.88877, 39.49435,
    28.24254, 25.05803, 33.45511, 37.8236, 22.1916, 17.92749, 18.77824,
    19.03162, 17.82331,
  91.94461, 105.2472, 107.033, 107.5656, 99.48592, 91.73083, 83.58383,
    77.19392, 60.36134, 51.47419, 62.72149, 65.0993, 72.28143, 72.84149,
    63.19975, 46.08965, 35.49227, 37.48937, 40.97271, 43.72961, 36.88481,
    29.3673, 36.37246, 31.03126, 24.34019, 19.63845, 18.31128, 18.11013,
    18.64655, 17.87722,
  82.19898, 87.52961, 89.39264, 85.81081, 75.6863, 76.70358, 91.92027,
    86.98054, 73.00756, 78.38235, 82.68631, 72.13023, 64.77991, 70.49775,
    67.79367, 47.95771, 45.03436, 46.80852, 51.21108, 51.03051, 40.17381,
    36.90289, 32.87065, 23.26488, 18.59204, 19.26429, 18.42097, 17.82418,
    17.71667, 17.28282,
  76.64931, 77.86718, 75.88033, 68.98576, 65.35329, 71.08473, 80.85671,
    75.69014, 69.04024, 70.32121, 68.60452, 57.20517, 50.60194, 57.34158,
    53.17603, 48.80257, 51.03617, 48.57713, 49.11884, 46.34618, 33.47543,
    28.18098, 23.30819, 20.47388, 19.79505, 19.11089, 18.35149, 17.9006,
    17.47803, 17.03556,
  66.5173, 62.92425, 56.1078, 53.08678, 54.31622, 56.09254, 61.29288,
    65.20609, 56.8463, 56.60752, 49.93517, 47.41101, 53.61764, 52.08768,
    50.04906, 49.94432, 48.77878, 43.46421, 43.42538, 40.72519, 25.00817,
    21.46671, 21.07739, 21.19067, 19.82133, 19.12443, 18.32754, 17.52662,
    17.3411, 17.06215,
  50.90328, 47.02686, 41.93472, 42.77628, 45.88663, 50.52333, 54.02906,
    53.96167, 49.15221, 44.04193, 43.75264, 52.91511, 57.11664, 56.73608,
    60.26978, 54.37914, 43.98366, 37.55973, 41.49548, 36.82283, 22.11509,
    22.41035, 22.30508, 21.41792, 18.98364, 18.70926, 18.31177, 17.15705,
    17.07659, 16.91431,
  44.67989, 41.75334, 37.10498, 37.17319, 41.89431, 45.6213, 44.72976,
    41.95577, 38.00204, 36.11009, 45.34957, 54.17027, 49.82317, 53.56334,
    54.3572, 45.85865, 42.32291, 43.01209, 45.35179, 38.50192, 27.14932,
    25.54506, 23.31423, 21.19874, 18.48583, 18.15824, 17.94304, 17.12093,
    16.95186, 16.82075,
  42.41721, 40.69906, 36.39315, 34.42199, 38.16287, 38.81115, 35.83577,
    33.21114, 32.43676, 40.48934, 50.24614, 47.13881, 44.3901, 46.30915,
    42.44733, 37.40208, 37.78974, 42.86084, 44.1288, 42.01526, 36.11881,
    29.70836, 23.55021, 21.17568, 19.09447, 18.17262, 17.74255, 17.22848,
    16.95024, 16.83789,
  39.8378, 39.6062, 34.63821, 32.52769, 34.04173, 33.3376, 30.7978, 29.87787,
    33.25138, 44.02665, 47.62664, 40.13626, 42.36766, 40.4193, 35.90145,
    33.43232, 34.31395, 37.20492, 38.73116, 38.90522, 35.77519, 31.53891,
    26.23829, 22.28728, 19.75802, 18.73615, 17.76099, 17.28714, 16.99627,
    16.85697,
  40.15128, 38.13742, 33.70559, 32.05188, 31.82272, 29.4006, 29.07892,
    30.53643, 37.14411, 44.89503, 41.79383, 36.31839, 38.26123, 35.09354,
    31.9584, 31.48039, 32.76083, 33.62774, 34.30101, 33.29281, 31.07088,
    29.59051, 27.44457, 26.54078, 23.14377, 19.84629, 18.01981, 17.47141,
    17.01377, 16.85252,
  38.98791, 37.51571, 32.23219, 30.07809, 31.12591, 31.6235, 32.38348,
    33.43362, 39.6488, 43.18766, 35.94802, 32.79152, 32.87947, 31.06131,
    29.81221, 31.69501, 33.38498, 31.89004, 30.18695, 28.34532, 27.51892,
    27.13859, 25.27538, 27.48756, 26.9391, 21.78524, 18.36645, 18.3077,
    17.53862, 16.9172,
  38.48996, 36.32627, 33.56863, 33.01641, 34.42009, 35.51427, 38.20454,
    39.47282, 43.75762, 41.22018, 31.97979, 31.16135, 31.59377, 31.84179,
    32.24741, 34.54755, 35.35624, 32.12753, 28.2514, 26.58839, 25.8201,
    24.91464, 24.24603, 25.32745, 26.30587, 24.7396, 21.40547, 19.14958,
    18.25503, 17.24009,
  36.8642, 38.60098, 33.18936, 32.64809, 35.67854, 37.41676, 38.96607,
    40.49419, 45.09889, 40.47992, 29.98586, 31.07793, 32.59951, 34.3718,
    35.90534, 37.43124, 35.43295, 31.88292, 27.47608, 24.35298, 24.57924,
    24.95409, 24.42257, 22.9845, 21.93354, 23.51237, 23.49772, 20.87649,
    19.95299, 18.3696,
  38.88197, 42.17327, 37.54921, 36.32916, 37.4248, 37.88341, 39.52533,
    42.7455, 43.96058, 36.89959, 30.36092, 32.4581, 35.23197, 36.90684,
    37.08293, 36.73114, 33.65186, 30.15728, 26.28478, 22.92839, 24.60966,
    25.94947, 23.17189, 20.32135, 19.45656, 21.18301, 23.64867, 22.62386,
    20.40332, 18.64138,
  42.2315, 45.33344, 41.34542, 38.77474, 38.74242, 37.69005, 40.75585,
    42.93295, 39.25405, 32.62223, 32.03135, 35.09575, 37.67104, 38.14393,
    36.7859, 34.51433, 31.24927, 28.1325, 24.92595, 22.48161, 24.49284,
    26.89162, 25.16899, 22.26572, 21.71796, 22.86617, 26.12597, 25.97035,
    20.34693, 17.4278,
  45.30986, 47.81979, 40.57584, 39.1673, 41.55563, 41.11433, 42.93494,
    41.18514, 33.40342, 31.30201, 33.75844, 36.91405, 38.47897, 38.01223,
    36.80707, 33.72995, 29.26076, 26.1877, 24.41059, 24.32231, 27.43757,
    29.12959, 26.56374, 24.20646, 23.51145, 24.57622, 26.33214, 28.95079,
    25.28795, 18.43814,
  40.64874, 36.59153, 37.33355, 42.71379, 45.52377, 48.00536, 45.68491,
    37.34597, 30.99339, 32.7434, 34.17067, 35.13628, 35.66504, 35.63477,
    35.44442, 33.11266, 29.75207, 28.21363, 26.15118, 25.08084, 26.9878,
    26.33767, 23.42807, 21.9213, 22.21266, 23.52243, 24.32527, 25.17445,
    24.87741, 20.07522,
  36.6528, 35.71042, 40.09935, 42.84344, 42.55763, 46.54719, 47.50472,
    36.6096, 30.96881, 34.13974, 35.61271, 36.78082, 37.40513, 37.34175,
    36.20738, 34.22242, 30.72409, 27.36696, 24.89236, 22.76996, 22.10919,
    21.2342, 20.38742, 20.07947, 20.63052, 21.76595, 22.39165, 21.3349,
    19.98802, 17.99946,
  19.45623, 19.78926, 20.14388, 20.59854, 20.80716, 21.10645, 21.54292,
    22.21234, 23.08863, 24.61673, 27.53709, 27.71132, 22.44801, 23.39461,
    23.76122, 22.46999, 22.89507, 24.36966, 26.27702, 29.43487, 31.49621,
    30.2008, 31.9245, 35.64784, 39.17875, 41.15103, 47.5927, 50.8326,
    29.39662, 22.89442,
  22.23492, 22.97656, 21.91682, 23.4597, 22.92761, 22.67103, 23.47855,
    24.22214, 25.25817, 26.63802, 28.66254, 30.92551, 31.8199, 28.80996,
    26.95337, 28.44367, 27.58083, 30.42925, 34.30051, 37.68555, 38.68958,
    39.42313, 42.57062, 50.55687, 58.20999, 55.1594, 49.41658, 52.95979,
    30.78704, 24.84586,
  20.22947, 20.4939, 20.78767, 21.24155, 21.49962, 21.98208, 22.52218,
    23.38096, 24.41303, 25.58543, 27.05483, 29.44674, 31.84064, 34.82953,
    37.2612, 36.00231, 39.21389, 43.87141, 47.52433, 53.41978, 62.0732,
    70.63933, 73.42799, 73.22196, 73.88521, 69.20832, 62.20307, 50.65435,
    31.46637, 26.94893,
  21.87948, 22.8373, 24.74372, 26.92822, 28.98213, 31.31032, 31.66585,
    31.22915, 32.46611, 34.48269, 35.51968, 36.74451, 38.68488, 40.82103,
    48.61312, 54.0715, 52.87637, 51.76177, 58.67247, 66.82431, 78.24871,
    81.29652, 74.72454, 80.54624, 80.88249, 77.85274, 69.73465, 49.58071,
    31.19069, 23.43512,
  26.94461, 26.35463, 29.27052, 31.26305, 32.8145, 32.51698, 32.14927,
    32.68398, 35.66995, 38.038, 37.41723, 39.43041, 43.03296, 48.36375,
    53.89204, 57.84005, 57.47392, 55.30699, 61.68656, 72.17556, 74.54945,
    62.26963, 63.23019, 71.42013, 78.06411, 76.86185, 67.88535, 71.53211,
    60.00331, 32.22312,
  28.16095, 30.9361, 35.11792, 39.38794, 38.36135, 35.70712, 37.51657,
    39.39627, 41.89192, 47.62226, 55.93739, 69.72621, 84.17104, 84.64412,
    88.30672, 94.05099, 95.08482, 84.43647, 72.2617, 71.41656, 63.27866,
    54.28939, 60.8362, 68.35023, 76.80984, 76.25336, 71.20778, 84.61983,
    71.47923, 30.24217,
  32.18056, 37.43193, 43.70346, 50.90859, 55.57007, 61.06808, 71.58638,
    83.14505, 86.27895, 86.7207, 87.34174, 81.27124, 72.03361, 73.4525,
    76.38981, 79.19518, 78.33436, 70.4821, 58.53578, 59.34761, 55.50549,
    55.043, 61.12946, 70.14568, 72.78844, 63.87769, 66.42873, 76.38889,
    59.72081, 22.17031,
  40.22849, 48.44727, 57.05305, 65.9942, 71.40327, 81.87794, 88.85597,
    73.10588, 62.30331, 61.8444, 56.37702, 50.83765, 46.39264, 48.17831,
    51.85409, 57.71655, 60.70499, 58.973, 51.25357, 52.12751, 51.7285,
    54.73616, 63.04991, 69.76822, 65.59169, 60.49503, 71.80438, 72.06095,
    46.7768, 22.91672,
  54.35556, 59.77193, 65.55078, 68.72393, 69.13919, 72.42469, 61.55315,
    54.49451, 55.84429, 55.28025, 53.85147, 53.68091, 58.38956, 73.05649,
    82.48918, 66.08288, 67.96069, 74.76699, 74.01685, 64.98071, 61.42355,
    74.84795, 88.72889, 88.13547, 72.53273, 78.20988, 77.64455, 62.08143,
    32.09639, 22.91146,
  79.57333, 88.91959, 85.73069, 88.60234, 79.54777, 67.91611, 48.45074,
    56.74662, 60.0416, 70.38365, 83.14764, 96.48224, 95.60735, 91.71949,
    84.3917, 92.3633, 98.37892, 96.54312, 88.1409, 84.15085, 91.82953,
    90.68137, 86.0322, 75.74004, 81.07671, 90.59649, 72.114, 39.70713,
    22.85954, 19.30832,
  102.0465, 96.46851, 95.61914, 86.35883, 97.59118, 98.61028, 94.70811,
    100.0131, 106.2554, 108.9695, 99.46474, 74.42184, 71.35728, 72.09908,
    76.31816, 84.11269, 89.05669, 87.15855, 82.27802, 80.82283, 90.34006,
    85.18, 64.38801, 55.6009, 61.73877, 60.9205, 39.36333, 22.69436,
    21.27209, 18.92608,
  104.0863, 90.92494, 103.601, 106.4212, 107.6134, 95.84898, 98.03572,
    90.57526, 80.20557, 68.25999, 60.90878, 57.0582, 64.61, 71.93053,
    75.67375, 76.82494, 74.7501, 72.02289, 67.46223, 67.80994, 75.48517,
    68.4185, 50.57665, 58.16579, 61.23421, 41.1858, 22.23017, 24.02208,
    22.35901, 20.07766,
  112.9318, 114.0553, 117.603, 118.0178, 116.3034, 111.1227, 95.51445,
    82.84882, 84.40947, 63.22404, 63.17611, 66.68854, 79.54445, 89.12627,
    84.95015, 71.23217, 71.32208, 66.60426, 62.6619, 68.5658, 71.24726,
    60.14013, 52.69984, 51.98272, 48.23076, 32.74455, 23.80919, 25.82431,
    24.76697, 21.94524,
  118.3706, 119.1174, 117.5316, 114.0154, 110.1182, 107.2552, 105.9859,
    105.4536, 101.8335, 101.9585, 103.6349, 102.3753, 105.3675, 106.881,
    104.3222, 87.04794, 85.73698, 89.83111, 93.83115, 88.52653, 71.98906,
    56.14688, 51.55264, 38.92755, 30.97083, 27.73084, 24.48562, 23.50928,
    23.32187, 21.69917,
  111.2638, 105.1838, 103.6656, 104.3506, 104.4725, 106.2019, 110.8268,
    110.6684, 106.6479, 107.0365, 106.0332, 105.1785, 106.5192, 106.659,
    105.4092, 105.0183, 105.0607, 103.8974, 101.5653, 87.39606, 55.81371,
    48.36744, 36.52296, 29.81993, 27.37653, 26.11991, 23.75582, 22.1427,
    21.07913, 20.06364,
  99.62182, 101.5808, 106.4083, 106.6763, 107.1171, 109.4927, 111.8314,
    108.8761, 106.4439, 106.1152, 106.2785, 104.013, 100.6725, 105.6616,
    104.922, 104.7766, 105.1287, 88.31215, 76.67765, 62.59174, 38.91032,
    37.12938, 30.39881, 28.57657, 27.25006, 24.98941, 22.81893, 21.77629,
    20.63838, 19.73823,
  89.81766, 89.20598, 92.84857, 97.44195, 101.7383, 105.7887, 106.7479,
    106.3185, 103.0834, 101.147, 94.09152, 104.2132, 107.3772, 105.4919,
    105.0566, 96.08643, 84.05269, 68.42079, 62.7798, 55.13803, 34.04045,
    34.9945, 30.9581, 28.67905, 26.35436, 25.08042, 22.63652, 20.63754,
    20.14582, 19.67503,
  74.31713, 78.80947, 79.17496, 83.17638, 86.01407, 90.09657, 91.88727,
    92.87982, 94.31646, 94.37758, 105.3607, 109.4579, 109.5811, 108.5658,
    108.2331, 90.47572, 66.39639, 56.08911, 61.35389, 54.00927, 34.94622,
    35.80064, 31.83099, 29.51816, 25.37516, 23.7719, 22.27674, 19.69158,
    19.57894, 19.25104,
  82.70993, 81.05705, 71.18566, 67.84018, 70.62878, 72.95348, 76.95541,
    82.50413, 87.07629, 97.24352, 107.413, 107.4793, 93.61094, 91.64803,
    84.85146, 75.33829, 74.55653, 77.20101, 79.6086, 66.75206, 45.49108,
    38.40025, 32.70127, 28.92792, 24.11403, 22.26695, 21.1988, 19.64421,
    19.31453, 19.14932,
  80.31374, 74.01401, 62.65511, 56.12674, 59.35974, 63.50672, 70.06757,
    77.48244, 86.96237, 100.3369, 102.6942, 80.80225, 71.93568, 69.76273,
    65.50113, 66.25082, 72.71013, 80.03743, 79.43993, 72.38391, 57.60993,
    43.53641, 33.38548, 29.11515, 25.56972, 22.48835, 21.19031, 19.9159,
    19.27923, 19.17574,
  70.37987, 63.3343, 54.03747, 50.29648, 54.75307, 60.77094, 67.15472,
    73.68623, 81.01916, 86.85193, 76.4494, 58.79727, 63.89937, 63.57125,
    62.78435, 62.96057, 66.18532, 66.79459, 65.09756, 59.97779, 53.2292,
    48.55632, 39.85271, 33.0666, 28.10616, 24.39935, 21.29413, 20.0896,
    19.31949, 19.2189,
  68.62098, 57.86415, 51.74173, 51.67223, 56.40518, 58.59525, 64.15827,
    67.52215, 73.38206, 73.60652, 59.4329, 51.61927, 58.7197, 59.80744,
    59.4291, 59.26242, 57.43151, 53.95797, 51.62528, 48.78488, 46.83729,
    45.35355, 43.48457, 41.83915, 34.77899, 25.95979, 21.73461, 20.54554,
    19.40893, 19.20126,
  63.47383, 57.13984, 51.78945, 52.63271, 61.42248, 65.67186, 66.11486,
    62.77693, 63.53679, 59.85075, 46.74823, 49.18513, 54.27121, 56.54305,
    55.16603, 55.03219, 52.73997, 46.01874, 43.02294, 42.16582, 41.78329,
    41.08601, 39.28646, 40.34131, 39.14875, 29.6822, 23.18073, 22.78714,
    20.82022, 19.32888,
  66.37487, 63.91637, 64.62955, 68.6273, 74.11694, 74.28221, 75.23236,
    70.38287, 69.10278, 57.56948, 45.91892, 53.61912, 58.3241, 60.83171,
    58.49183, 56.3243, 53.7159, 47.8212, 42.29523, 40.75904, 39.57093,
    37.95123, 36.20486, 35.6218, 36.42468, 35.50419, 29.95736, 24.46018,
    22.51786, 20.21453,
  70.39108, 73.65321, 69.48297, 71.69663, 75.40328, 73.9163, 70.10921,
    68.83285, 71.93028, 61.31889, 48.66139, 57.55843, 60.93753, 62.56927,
    59.99036, 58.31094, 53.31872, 48.52274, 43.67307, 39.27611, 38.63851,
    38.21673, 35.41968, 32.66069, 32.35605, 35.85389, 36.48572, 30.49999,
    26.71423, 23.07219,
  83.2326, 87.45587, 84.1954, 79.8355, 75.42168, 71.74646, 74.21985,
    77.24766, 71.03088, 58.73005, 55.49224, 61.84481, 64.0589, 61.59098,
    56.71294, 54.80378, 51.81933, 48.20636, 45.21313, 40.61187, 39.42292,
    38.16777, 33.65523, 30.7783, 31.94414, 35.26033, 38.32076, 34.48212,
    26.7954, 22.83211,
  94.05284, 94.44984, 83.87193, 76.45383, 72.62894, 69.04619, 76.22173,
    76.2812, 63.77333, 55.84023, 60.91555, 64.3661, 63.10082, 59.15217,
    55.39259, 52.65334, 49.74307, 46.51297, 42.90911, 39.30737, 40.33662,
    43.66114, 43.05522, 39.8829, 40.0817, 42.01941, 45.36261, 41.48877,
    27.19643, 20.22792,
  97.30058, 90.61652, 80.79236, 78.74667, 78.8694, 76.90123, 78.84082,
    71.75774, 57.98954, 59.92039, 62.91312, 63.07195, 60.86971, 58.13862,
    56.19587, 52.50845, 47.40492, 45.3038, 46.15371, 48.42854, 50.79094,
    50.46313, 46.87531, 45.00464, 44.85203, 46.65605, 47.72277, 48.9548,
    40.10027, 23.70729,
  82.71616, 77.40543, 80.88569, 89.91978, 89.76121, 90.71906, 82.00041,
    64.84381, 56.90398, 58.60198, 54.16785, 51.3129, 51.25977, 52.66167,
    54.73271, 54.63412, 53.74807, 54.68301, 53.33862, 50.24288, 49.53634,
    46.32711, 42.6158, 40.91205, 41.72337, 42.78478, 42.17124, 39.22265,
    35.48694, 27.09651,
  81.03621, 83.15572, 85.17123, 84.09708, 84.68874, 90.83696, 88.06625,
    66.04097, 55.22179, 58.00034, 58.2859, 60.74567, 63.04922, 64.27885,
    63.31896, 61.09253, 55.73919, 49.33783, 46.21707, 42.51198, 39.41246,
    37.63255, 36.27991, 35.36044, 35.10408, 35.07868, 33.73844, 29.32853,
    25.00481, 20.47653,
  26.16023, 26.52771, 27.08319, 27.82772, 28.4809, 29.41481, 30.5438,
    31.90223, 33.52006, 35.68566, 38.90034, 40.02109, 37.22698, 38.69299,
    39.7182, 39.32726, 39.87664, 41.1694, 42.71651, 44.96505, 46.11411,
    44.78916, 45.57214, 47.96635, 49.65329, 49.43242, 52.97276, 53.98281,
    38.07833, 32.6167,
  27.54152, 28.42085, 28.42083, 30.39617, 31.09298, 32.26497, 34.34319,
    36.48207, 38.89144, 41.69119, 45.17313, 48.94997, 51.25909, 50.03752,
    49.43878, 50.44785, 49.71041, 51.26141, 53.40353, 55.30751, 55.66142,
    55.19506, 55.3942, 58.41945, 61.90519, 57.33311, 50.05964, 53.15495,
    38.70018, 34.03875,
  29.1151, 30.83985, 32.63845, 34.62162, 36.59378, 38.6415, 40.65587,
    42.86795, 45.18142, 47.55544, 49.9843, 52.82121, 55.38402, 58.13119,
    59.70884, 57.77271, 59.27709, 61.94172, 64.54488, 69.05154, 75.73351,
    81.13374, 80.25481, 75.74585, 72.87691, 69.1409, 61.35006, 50.67104,
    37.92128, 34.76321,
  36.29366, 39.11586, 42.45258, 45.81647, 48.72859, 51.49102, 52.70199,
    53.22378, 54.65075, 56.2364, 56.88688, 57.48142, 57.56529, 57.44188,
    61.46538, 63.68273, 61.11024, 59.9565, 65.1891, 71.2505, 79.76942,
    80.86656, 75.47167, 79.89066, 78.50752, 76.58264, 72.13351, 56.34745,
    40.81385, 33.26511,
  44.37623, 46.64527, 50.83888, 54.01874, 56.36741, 57.65251, 58.77216,
    59.88157, 62.54411, 64.50122, 64.71771, 67.18162, 68.73622, 69.0163,
    69.87858, 70.51952, 67.47649, 63.09194, 65.51517, 72.28966, 73.08501,
    64.32043, 66.66213, 73.40332, 79.67946, 80.27731, 75.12964, 79.21771,
    68.33228, 42.05165,
  58.37778, 64.57317, 69.77911, 74.63124, 74.74556, 74.44408, 77.23405,
    77.45956, 77.27333, 79.61786, 84.34907, 93.8876, 102.9518, 99.41536,
    98.79428, 99.22246, 95.43472, 85.40407, 74.16409, 71.30917, 64.03703,
    56.87875, 62.43644, 67.40311, 73.08125, 73.02457, 71.69139, 84.01785,
    73.69643, 37.49384,
  67.19284, 72.15393, 76.39835, 80.55328, 82.33424, 85.18726, 90.94556,
    94.82237, 92.29809, 87.49385, 83.62063, 73.76933, 62.6524, 64.44656,
    66.4749, 69.29417, 70.51147, 66.61226, 59.79762, 61.05729, 58.88615,
    58.43598, 62.48219, 68.35567, 69.46891, 64.81741, 68.31095, 75.23959,
    60.84759, 31.06233,
  60.86512, 64.70409, 69.43438, 73.90895, 76.25319, 83.49054, 85.42596,
    68.57127, 60.79266, 62.01476, 59.93723, 58.17305, 57.55964, 60.1382,
    62.48285, 65.8953, 69.05759, 67.60144, 62.23597, 62.66095, 63.68837,
    66.4862, 71.23924, 73.78479, 69.89499, 68.68179, 76.10872, 73.38304,
    51.28513, 32.65911,
  70.31305, 73.54409, 77.49153, 80.26676, 82.05032, 85.30465, 77.92162,
    79.0916, 83.64024, 85.98927, 87.48298, 88.28307, 90.92966, 99.65993,
    102.3565, 88.92786, 87.18085, 88.58154, 85.19212, 77.60437, 74.48758,
    81.34677, 87.76625, 84.60136, 74.40062, 78.49142, 76.535, 61.48033,
    36.40565, 32.57151,
  98.97946, 105.8001, 98.56984, 99.88088, 100.7936, 94.8767, 78.93533,
    88.01497, 89.00844, 93.33107, 98.94129, 105.7276, 102.6939, 97.27464,
    91.98134, 96.25008, 97.5857, 93.65822, 88.19941, 86.92456, 88.99316,
    84.01912, 77.19547, 68.32238, 72.28752, 79.26033, 67.03706, 43.22572,
    31.84667, 29.83092,
  111.0486, 110.5625, 112.3632, 107.5506, 114.4675, 108.5662, 99.54439,
    101.0029, 100.366, 93.58876, 79.92811, 63.50987, 60.8832, 61.49911,
    62.32504, 64.34772, 67.30468, 68.23102, 68.6856, 71.94191, 80.99648,
    75.37141, 60.84045, 57.67705, 62.31135, 58.4596, 42.01018, 32.53851,
    32.2371, 29.96125,
  115.8235, 112.193, 115.333, 116.4295, 116.9604, 101.1978, 97.30747,
    87.78633, 77.92521, 67.42122, 62.24606, 59.41711, 62.24018, 63.23702,
    61.0149, 59.73072, 58.52012, 58.85347, 59.77752, 64.627, 72.56828,
    70.33154, 59.88688, 67.37928, 68.95838, 52.26206, 33.93042, 37.55902,
    33.72302, 31.32188,
  123.4582, 123.5537, 125.534, 126.6918, 126.287, 122.7493, 115.3331,
    105.668, 110.0719, 91.99884, 86.91843, 81.98796, 88.37616, 90.42151,
    80.08082, 65.40917, 66.66285, 64.92109, 64.10176, 68.75077, 70.28939,
    63.75837, 57.23277, 53.14146, 51.748, 44.54785, 35.63736, 36.97582,
    35.95776, 32.76401,
  112.1994, 112.7421, 113.1821, 113.6549, 114.0133, 114.8326, 116.0055,
    117.112, 115.7259, 116.4281, 117.8104, 116.6817, 118.0366, 118.5162,
    106.2598, 84.93875, 80.11942, 83.20061, 84.61626, 75.81721, 63.72234,
    54.07083, 48.79218, 40.76819, 36.55606, 35.73994, 33.43579, 32.62813,
    32.99792, 32.02018,
  107.0749, 104.1363, 109.0609, 111.2563, 112.5989, 114.4068, 116.8691,
    117.1683, 114.3392, 111.7878, 103.2903, 95.51051, 96.31006, 97.87358,
    96.2887, 92.38502, 81.54723, 76.84508, 75.54698, 67.79423, 49.92022,
    48.63315, 41.12532, 38.22739, 37.16911, 35.35484, 33.60197, 32.29181,
    31.21896, 30.54139,
  107.7168, 111.4316, 112.2396, 112.4848, 111.774, 113.5962, 114.4942,
    104.4145, 91.98057, 85.3709, 82.29485, 75.42041, 70.95256, 78.05447,
    75.39225, 73.63607, 73.70187, 64.40042, 61.29103, 54.58339, 42.61406,
    44.22234, 39.73656, 38.23592, 37.23343, 35.20538, 33.22027, 32.40846,
    31.45625, 30.60575,
  90.36945, 89.09261, 91.00886, 93.51616, 95.48438, 97.39794, 97.41649,
    95.61923, 91.49139, 84.17554, 75.60735, 83.15172, 90.96866, 81.33713,
    74.44116, 68.95997, 63.57331, 59.46796, 59.31015, 54.73552, 43.29409,
    44.68464, 40.87247, 38.3459, 36.53796, 35.35343, 32.81376, 30.94197,
    30.79324, 30.45944,
  81.15587, 85.1233, 84.9792, 87.73395, 89.36911, 91.24591, 90.68545,
    90.09113, 89.18232, 87.76826, 96.07718, 104.1466, 99.47745, 95.00338,
    88.17345, 76.35045, 67.10412, 63.95742, 66.24772, 58.63241, 44.52425,
    43.9702, 41.13111, 39.31081, 35.76906, 33.97595, 32.78606, 30.30524,
    30.27726, 30.05413,
  92.67924, 86.68492, 75.29533, 68.86476, 69.02345, 68.11173, 69.2581,
    70.44518, 71.52721, 76.24913, 83.87367, 82.6033, 73.77608, 77.51909,
    79.54541, 81.57943, 88.76582, 93.62784, 89.96125, 77.07132, 57.01085,
    47.7051, 42.45656, 39.45731, 35.52523, 33.36805, 32.22721, 30.67915,
    30.19314, 30.0762,
  87.47882, 78.09223, 65.18877, 57.8464, 58.70024, 60.31063, 62.78299,
    65.73318, 69.87753, 76.03444, 76.12134, 64.37965, 64.07841, 63.77273,
    62.58408, 63.28913, 68.58273, 74.99004, 77.31092, 75.3445, 66.61877,
    55.6645, 46.55509, 42.47009, 38.73333, 34.48524, 32.56961, 30.92549,
    30.16771, 30.08695,
  78.68568, 69.69881, 60.12732, 53.39422, 55.59169, 57.65617, 59.73583,
    61.20967, 63.37065, 65.4019, 58.8161, 50.41162, 54.42146, 53.61814,
    52.24843, 51.24683, 53.40156, 56.15678, 59.84806, 61.5645, 61.9537,
    61.82786, 55.10826, 47.6453, 41.41447, 35.95455, 32.55796, 31.05956,
    30.16931, 30.08471,
  76.74162, 68.5202, 59.28571, 57.11292, 57.85662, 56.40906, 56.92144,
    56.111, 58.37977, 57.25914, 47.67337, 42.64309, 45.8343, 45.83243,
    44.84945, 45.35187, 45.59068, 46.90903, 49.96297, 52.00031, 53.03517,
    53.64973, 54.64258, 53.66004, 46.7743, 37.39159, 33.36995, 31.99877,
    30.42859, 30.0466,
  77.57768, 73.24666, 65.95107, 62.58739, 66.40287, 65.08494, 61.53951,
    56.25589, 55.47868, 51.86848, 43.51929, 45.48868, 46.97479, 47.73124,
    46.8175, 47.89418, 47.95695, 45.5029, 45.67561, 46.85253, 47.67466,
    48.01285, 47.86613, 50.27418, 50.9762, 42.79417, 36.02587, 34.4747,
    32.1749, 30.22464,
  86.88678, 85.2422, 80.94568, 79.54795, 78.79984, 76.58637, 76.52439,
    73.84354, 73.67641, 65.37101, 57.1696, 61.20234, 62.71425, 63.52862,
    61.17669, 59.54957, 58.04533, 54.75274, 51.21461, 50.41565, 49.67965,
    48.83121, 48.03822, 47.93383, 50.16323, 50.60068, 44.58299, 37.5827,
    34.80584, 31.50206,
  85.19212, 82.12657, 73.79685, 71.41811, 71.85378, 71.25645, 71.50062,
    75.11494, 79.08447, 69.76912, 59.88565, 63.82415, 65.70618, 66.53852,
    64.99461, 64.01505, 61.01547, 58.8059, 56.73178, 54.14905, 52.81846,
    51.2807, 48.14943, 46.59117, 48.18153, 51.58829, 52.03901, 43.94109,
    37.87597, 33.78426,
  94.65759, 90.80137, 83.02941, 76.55138, 73.07639, 72.75172, 77.40681,
    80.62904, 75.76115, 66.30322, 64.30572, 66.18774, 67.79626, 66.69547,
    63.87132, 63.30293, 62.1521, 61.00487, 61.07324, 59.32116, 57.8924,
    56.08167, 51.93064, 49.15957, 50.03209, 51.79959, 53.44363, 46.4854,
    36.18952, 32.7815,
  96.25626, 89.49778, 79.31636, 73.6495, 71.29647, 68.3289, 73.6055,
    73.44327, 66.73413, 62.73841, 66.37997, 68.64386, 69.86902, 69.43755,
    68.3677, 67.10113, 65.55965, 65.45369, 65.88561, 65.79215, 66.39059,
    67.54287, 65.72988, 62.07021, 61.59858, 62.46205, 63.81926, 56.80074,
    39.60543, 30.97926,
  95.61041, 88.37496, 83.3951, 81.23535, 79.71282, 75.9381, 73.57361,
    68.66067, 61.66349, 64.16428, 66.82709, 69.58128, 71.30653, 72.05529,
    72.27374, 69.98604, 66.4574, 65.71206, 67.0433, 67.75577, 65.16293,
    60.2972, 56.55818, 55.35291, 56.36219, 57.97071, 59.05046, 60.54425,
    51.97286, 35.13518,
  81.64034, 77.96713, 79.9025, 82.2468, 83.8634, 85.30208, 77.1082, 64.36979,
    60.18564, 61.3042, 59.37627, 58.68714, 59.31139, 60.02599, 60.46282,
    59.33791, 56.65899, 54.885, 51.93615, 48.66821, 47.57518, 45.71174,
    42.94317, 41.22343, 42.19637, 43.41785, 43.46907, 41.64985, 40.99649,
    36.34466,
  73.94583, 73.61494, 72.36232, 71.35156, 76.33449, 84.35942, 84.13504,
    68.33987, 61.53506, 64.38396, 64.85384, 64.84048, 63.6498, 60.66547,
    55.73483, 51.2341, 44.93668, 39.95333, 39.50406, 38.62832, 36.97026,
    37.1876, 37.1498, 36.9888, 37.3679, 38.44713, 38.54591, 35.72582,
    32.4009, 30.06845,
  38.24385, 39.228, 39.90129, 40.68124, 41.29617, 42.0322, 42.76532,
    43.51832, 44.3457, 45.40322, 46.91891, 46.98123, 44.52167, 44.67916,
    44.5465, 43.53011, 43.26721, 43.46482, 43.88012, 44.8139, 44.94669,
    43.45408, 43.91595, 45.89509, 47.33951, 46.69886, 48.71104, 50.0703,
    38.94454, 34.93098,
  44.25359, 45.5101, 45.61993, 46.91125, 47.19184, 47.79211, 48.91208,
    49.95134, 51.11672, 52.36422, 53.88027, 55.48767, 56.09382, 54.51937,
    53.33408, 53.28607, 52.26101, 52.7267, 53.59001, 54.36053, 53.99597,
    53.08593, 53.06882, 55.78703, 58.35962, 52.85595, 45.83938, 48.3026,
    39.2343, 35.71656,
  47.42923, 48.64574, 49.31162, 49.95514, 50.44944, 51.13634, 51.88585,
    52.75747, 53.69189, 54.59274, 55.52757, 56.77758, 57.88031, 59.30374,
    60.03458, 58.38038, 58.93457, 60.54359, 62.27245, 65.26619, 70.24068,
    74.63565, 74.07739, 70.48297, 67.5515, 62.25443, 55.13117, 46.59311,
    38.44695, 36.3262,
  52.97107, 54.33118, 55.54854, 56.64214, 57.31204, 58.17709, 58.36713,
    58.14416, 58.56487, 59.04776, 59.07851, 59.02446, 58.50671, 57.70975,
    59.79566, 60.70773, 58.52173, 57.62648, 61.03004, 65.09992, 71.22334,
    71.67111, 67.17043, 70.45449, 68.20874, 66.6557, 63.22986, 52.274,
    40.61234, 35.38717,
  60.26599, 60.76762, 62.02419, 62.68313, 62.73258, 62.59283, 62.99484,
    63.19149, 64.42767, 65.24912, 65.41302, 67.24854, 67.73259, 66.48303,
    66.3261, 66.41347, 63.7831, 60.06551, 60.45023, 64.59398, 64.26033,
    56.73411, 58.12045, 63.19545, 67.31915, 67.08104, 64.66385, 69.80168,
    63.88441, 42.52484,
  65.11066, 67.8343, 70.214, 72.34302, 71.33866, 70.8524, 73.45382, 73.93667,
    73.13414, 73.75505, 76.71304, 84.4433, 91.5818, 87.83669, 87.07312,
    88.07961, 85.5598, 77.5674, 68.25716, 64.6811, 57.67568, 51.07189,
    55.2241, 58.78098, 62.95248, 63.61559, 64.61731, 74.92258, 66.29043,
    39.15701,
  65.69577, 69.39262, 72.42471, 75.3568, 76.7589, 79.49223, 85.64264,
    90.51164, 88.64402, 83.63589, 79.66725, 71.08753, 61.14171, 61.53856,
    61.91911, 63.20963, 63.85545, 60.52795, 55.61613, 55.79602, 53.31744,
    52.32407, 55.0164, 58.85804, 59.8755, 57.62303, 60.49455, 66.53024,
    56.31944, 33.66497,
  70.35977, 74.0752, 77.22195, 80.22629, 81.71659, 86.87721, 88.72369,
    75.76471, 69.26019, 68.95966, 66.0724, 62.99229, 60.78462, 60.33525,
    59.97144, 60.64383, 62.03209, 60.62706, 56.77409, 56.30316, 56.23417,
    57.76162, 60.81451, 62.50219, 60.20798, 60.0351, 65.66965, 64.05434,
    47.44006, 34.38223,
  80.14247, 81.3191, 82.14537, 83.09911, 84.39647, 85.08957, 76.9613,
    76.15547, 78.54668, 78.56156, 78.23582, 77.38749, 77.47733, 82.08812,
    83.04486, 73.97868, 72.92458, 73.14018, 70.58295, 64.93728, 62.12383,
    65.74751, 70.05715, 68.36787, 62.97843, 67.05563, 67.29333, 55.77325,
    36.66105, 34.64066,
  92.16992, 93.41161, 86.32091, 85.77946, 86.61803, 80.43902, 65.86073,
    71.00193, 70.23505, 71.72778, 73.98753, 77.87227, 76.56348, 73.93369,
    71.9964, 76.03461, 77.55893, 75.05418, 71.79818, 70.71149, 71.35625,
    67.68871, 63.17996, 57.2923, 60.88444, 67.87275, 60.807, 42.37183,
    34.10145, 33.09277,
  114.3672, 113.5831, 107.9595, 95.10445, 96.24211, 87.30879, 78.18262,
    78.38615, 78.04497, 74.05803, 64.35294, 53.98746, 52.94606, 53.69354,
    54.83073, 56.58886, 58.45723, 58.94096, 59.49303, 61.78799, 67.43048,
    64.24809, 54.91154, 53.14609, 56.49908, 53.981, 42.0398, 34.29687,
    34.52795, 33.13474,
  123.4046, 120.4102, 121.4774, 120.3138, 117.2287, 96.51278, 89.90178,
    80.70135, 73.44962, 67.18013, 62.599, 59.45515, 60.91608, 60.33141,
    56.68912, 55.51571, 54.28865, 53.81939, 53.91392, 56.79292, 61.80706,
    60.61205, 54.61499, 60.07674, 61.67378, 48.91914, 35.29077, 37.92737,
    35.33617, 33.93266,
  126.1096, 126.6725, 127.3583, 126.5974, 124.1377, 119.6811, 112.0758,
    100.6747, 102.6868, 89.23228, 83.4214, 77.8091, 81.21562, 81.901,
    72.55775, 59.66612, 60.35643, 59.0426, 57.52444, 59.26594, 60.21083,
    56.84248, 52.54872, 48.27625, 47.42138, 42.79364, 36.6798, 37.62675,
    36.97065, 34.91963,
  112.956, 113.3057, 109.5357, 107.497, 106.0182, 110.8823, 113.2361,
    112.4785, 101.0941, 102.7179, 105.5561, 99.48529, 98.42781, 96.69727,
    87.98141, 73.5349, 67.91479, 71.67097, 72.80611, 66.14465, 57.91883,
    51.21572, 45.85861, 39.87026, 36.72754, 36.7919, 35.60987, 34.9252,
    35.20789, 34.49405,
  78.84947, 75.11431, 77.08128, 77.92984, 79.45612, 82.07417, 86.71708,
    84.11769, 80.14726, 79.88812, 76.60274, 72.94615, 75.15688, 78.42574,
    77.74454, 75.15092, 69.35971, 65.57844, 64.27998, 59.08526, 47.41869,
    46.11655, 40.83387, 37.9309, 37.69621, 36.83378, 35.74959, 34.71167,
    33.96646, 33.50605,
  76.66682, 78.51979, 78.77755, 78.15189, 77.70899, 79.63989, 81.50353,
    76.44784, 70.05891, 66.86537, 65.88739, 62.38283, 60.90063, 64.82517,
    62.90703, 62.15208, 62.79107, 57.00658, 54.13772, 49.31592, 42.03163,
    42.3773, 39.13967, 38.07199, 37.62633, 36.77859, 35.5551, 34.83389,
    34.16207, 33.54318,
  68.70409, 67.74049, 68.52309, 70.22873, 71.91762, 73.59512, 75.44513,
    76.79964, 74.90565, 71.32481, 66.52194, 70.9718, 75.29125, 69.8563,
    64.06094, 60.35387, 57.00956, 53.95448, 52.81148, 49.41916, 42.13338,
    42.47482, 39.63023, 38.0374, 37.24856, 36.77608, 35.13261, 33.84447,
    33.66468, 33.42825,
  64.56267, 65.43339, 64.43192, 66.53415, 68.7388, 71.39359, 73.39775,
    75.30815, 76.16311, 75.30226, 79.84383, 83.50384, 81.27657, 79.45026,
    75.23843, 68.99513, 63.88633, 61.44809, 60.6291, 54.07328, 44.05873,
    42.31033, 40.08621, 38.84823, 36.88144, 35.77884, 34.89689, 33.39362,
    33.3143, 33.16864,
  72.63942, 67.44048, 59.56803, 56.48864, 58.78329, 59.59616, 61.31245,
    62.8657, 63.02694, 65.21738, 68.92398, 67.55336, 62.90826, 65.44111,
    66.39158, 68.78571, 74.74497, 78.46761, 75.76289, 66.6692, 53.48157,
    45.62807, 41.53439, 39.6382, 37.16637, 35.60393, 34.67299, 33.60262,
    33.24901, 33.15402,
  66.06979, 60.79073, 53.2923, 49.05888, 50.88763, 51.92232, 53.37189,
    54.86237, 56.97286, 60.91346, 60.99266, 54.81972, 54.85311, 54.09918,
    53.36426, 54.23572, 58.15443, 63.23937, 65.04196, 63.82423, 58.26178,
    50.71886, 44.37056, 41.64478, 39.27597, 36.49495, 34.99693, 33.72959,
    33.21569, 33.17141,
  60.45294, 56.02068, 48.8699, 45.25187, 46.26283, 47.12552, 48.48092,
    49.98739, 52.30645, 54.5799, 51.85592, 48.07449, 50.82838, 50.08422,
    48.55949, 48.22285, 49.57829, 51.35118, 53.21056, 53.20127, 53.1656,
    53.03011, 49.13182, 44.98535, 41.15896, 37.48726, 34.98769, 33.86357,
    33.22955, 33.19061,
  63.07064, 59.65846, 52.85448, 50.09542, 50.53002, 49.15508, 49.72317,
    50.24917, 52.77293, 53.04395, 48.16965, 45.71967, 47.29486, 47.03014,
    46.20499, 46.30119, 45.99848, 46.28931, 47.57483, 48.21534, 48.0154,
    47.84208, 48.58984, 47.86477, 43.96872, 38.35439, 35.49191, 34.44026,
    33.41305, 33.18239,
  70.06455, 69.48192, 62.58571, 60.44341, 62.52128, 62.16061, 60.16627,
    57.52621, 57.61805, 55.81951, 51.08363, 51.38593, 51.6258, 51.37391,
    49.92122, 49.72432, 48.93048, 46.76936, 46.12149, 45.95621, 45.51871,
    44.85076, 44.32729, 45.64692, 46.18378, 41.6106, 37.26989, 36.03891,
    34.48162, 33.28428,
  76.23491, 75.89629, 72.01031, 70.81879, 70.55836, 69.21236, 69.84803,
    69.6162, 70.75427, 66.12544, 61.39202, 63.26727, 64.21346, 63.98658,
    61.46855, 59.23953, 56.9119, 53.73812, 50.7305, 49.23495, 47.58106,
    46.15541, 45.30308, 44.9445, 46.30624, 46.68124, 42.92667, 38.11965,
    36.23346, 34.13365,
  78.16092, 74.77261, 68.49066, 66.75593, 66.99612, 66.33992, 67.78868,
    71.44384, 74.99567, 69.67886, 63.18544, 65.16835, 65.7801, 65.59452,
    63.63199, 61.72084, 58.34184, 55.83998, 54.0012, 51.70195, 49.92362,
    47.94012, 45.58347, 44.28504, 45.32738, 47.53104, 47.4866, 41.83961,
    38.00459, 35.48944,
  83.71445, 81.5808, 76.08079, 70.90816, 68.92026, 68.60187, 72.72418,
    77.26637, 75.86261, 69.48415, 68.0268, 68.43285, 68.81921, 67.29424,
    64.40385, 62.57466, 60.26945, 58.17966, 57.28993, 55.59155, 54.13842,
    52.17123, 48.67654, 46.23814, 46.40432, 47.12363, 47.81186, 43.14945,
    36.83987, 34.77889,
  85.41874, 82.46009, 75.45091, 71.35049, 68.4117, 66.28854, 69.89483,
    71.32669, 68.65553, 65.99342, 67.3201, 68.04357, 68.22685, 67.52349,
    65.60497, 63.53947, 61.62352, 60.36037, 59.79248, 58.82877, 58.43981,
    58.46925, 56.64532, 53.74989, 52.84256, 53.11781, 54.01346, 49.5132,
    38.91326, 33.70554,
  79.75416, 77.39247, 73.80035, 72.39334, 70.55012, 67.03329, 64.85276,
    61.71262, 57.68908, 58.02281, 58.58303, 59.89702, 61.18911, 61.77278,
    61.61681, 60.19683, 57.94089, 57.06009, 57.6233, 57.76343, 56.05039,
    53.13863, 50.54373, 49.38139, 49.70272, 50.55067, 51.14701, 52.0273,
    46.67434, 36.31703,
  61.82272, 60.68711, 61.85903, 62.93894, 64.69464, 66.07336, 60.74995,
    52.27254, 49.64052, 50.36668, 49.42611, 49.35221, 50.0873, 50.52508,
    50.59843, 50.49769, 49.50678, 48.76159, 47.26442, 45.43686, 44.74549,
    44.0186, 42.56639, 41.30472, 41.70335, 42.10251, 41.7155, 40.57788,
    40.15877, 37.06636,
  50.04566, 50.19576, 49.51129, 48.52263, 50.8005, 55.49459, 56.00679,
    48.11581, 44.74782, 47.26607, 48.72833, 49.9594, 50.34478, 48.96912,
    46.55368, 45.07447, 41.99749, 39.33671, 39.05711, 38.56892, 37.62684,
    38.09404, 38.42227, 38.31156, 38.34462, 38.79142, 38.52844, 36.83537,
    34.8762, 33.28009,
  38.64885, 38.81541, 38.98822, 39.14844, 39.22173, 39.42736, 39.68038,
    40.0063, 40.44152, 41.16137, 42.29126, 42.31845, 40.59346, 41.12081,
    41.3177, 40.85418, 41.20615, 41.91632, 42.75551, 43.95248, 44.37615,
    43.42681, 44.08758, 45.85812, 47.35999, 47.49178, 49.17926, 49.90408,
    41.72254, 38.98217,
  42.57865, 42.85237, 42.32765, 42.82245, 42.56158, 42.54122, 42.88248,
    43.17073, 43.5721, 44.17565, 44.97828, 46.01702, 46.61576, 45.56243,
    44.87475, 45.44879, 45.23532, 46.41073, 47.84424, 49.017, 49.25794,
    49.32669, 50.59669, 53.94597, 56.87724, 52.78959, 46.54544, 49.28241,
    42.24131, 39.68054,
  45.56573, 45.89355, 45.97793, 46.14371, 46.29696, 46.5884, 46.96205,
    47.4789, 48.03519, 48.6408, 49.42265, 50.59523, 51.72391, 52.9403,
    53.67191, 53.01464, 54.31519, 56.3673, 58.33018, 61.24984, 65.72321,
    70.2027, 70.35577, 66.62937, 63.84251, 59.87813, 54.22773, 48.09174,
    42.00294, 40.30224,
  49.6568, 50.26627, 50.96881, 51.756, 52.41471, 53.24889, 53.52292,
    53.54527, 53.99728, 54.54288, 54.93648, 55.60201, 55.78862, 55.38152,
    57.41001, 58.80315, 57.75391, 57.57628, 60.72008, 64.26511, 69.4169,
    69.11559, 63.41368, 65.2225, 62.98731, 61.27959, 59.57171, 50.39132,
    42.12183, 39.26193,
  52.69354, 52.40251, 53.14895, 53.59733, 53.78419, 53.87643, 54.47234,
    54.89909, 55.89233, 56.46772, 56.41566, 57.81859, 58.80408, 59.06734,
    60.04844, 61.37936, 60.51673, 59.09265, 61.28052, 65.60925, 65.23694,
    57.58911, 57.30983, 60.75036, 63.77396, 64.17524, 62.13924, 66.57079,
    62.56438, 46.39679,
  59.05395, 61.14368, 63.17513, 65.16485, 64.83277, 65.08956, 67.78864,
    68.94746, 69.78736, 71.69164, 75.42076, 83.69846, 91.01115, 88.0316,
    87.86537, 88.78311, 86.47575, 79.58192, 71.19394, 67.63772, 61.00761,
    54.95996, 58.56342, 61.28352, 64.83096, 65.5759, 66.4638, 75.90796,
    69.84076, 43.46404,
  64.94453, 67.80077, 70.25034, 72.78401, 74.16483, 77.196, 83.76724,
    88.9313, 87.95163, 83.94711, 80.18714, 72.6724, 64.01466, 64.60957,
    65.13332, 66.38089, 66.78069, 63.49223, 58.94833, 57.92585, 55.11517,
    54.3385, 56.87005, 60.34513, 61.69855, 60.34708, 64.13999, 69.96342,
    59.09861, 38.10626,
  63.1594, 65.18322, 67.24873, 69.20528, 70.11432, 74.79842, 76.57797,
    64.02477, 57.54146, 57.40208, 55.10715, 52.8869, 51.68646, 52.53886,
    53.6791, 55.89111, 58.149, 57.81525, 55.35722, 55.26934, 55.32419,
    56.75452, 59.78504, 62.27299, 61.71662, 62.875, 68.88528, 67.03061,
    51.4782, 38.38468,
  67.49261, 68.4993, 69.63811, 70.39422, 71.86522, 72.58611, 64.61395,
    62.79688, 64.66955, 64.69135, 64.88814, 65.16498, 66.60583, 71.34245,
    73.13316, 66.92977, 67.2325, 68.96825, 67.90056, 63.87855, 62.16508,
    65.46173, 69.12811, 68.15845, 65.0224, 69.81859, 70.54592, 59.36948,
    40.63125, 38.93234,
  77.20302, 80.4758, 76.01071, 76.88039, 79.03773, 74.48604, 62.13012,
    67.21496, 67.45851, 69.6123, 72.11202, 76.08719, 75.74142, 73.99087,
    72.14059, 74.58317, 75.5682, 74.29386, 72.47388, 71.35735, 71.70311,
    69.19679, 65.74888, 61.40626, 65.50697, 72.11159, 64.40952, 46.19072,
    38.24947, 37.68979,
  100.7446, 97.38091, 92.78878, 82.79247, 85.57203, 78.83845, 71.45238,
    73.50034, 74.1299, 71.42471, 63.89217, 55.45754, 55.26764, 56.17964,
    56.92756, 58.33527, 59.92315, 60.44617, 60.85233, 62.68011, 67.06844,
    64.44945, 56.99469, 55.77972, 59.94421, 58.22556, 46.49633, 38.19442,
    38.63675, 37.65518,
  106.9203, 103.9115, 105.5584, 105.4379, 97.98738, 80.35472, 77.39459,
    69.99361, 63.58241, 60.12899, 56.63318, 55.09959, 56.94617, 56.85336,
    55.12133, 55.0707, 54.75342, 55.15044, 55.6664, 58.09811, 62.77961,
    62.2647, 57.53849, 62.83215, 64.11417, 51.91828, 39.00492, 41.10909,
    39.05001, 38.19301,
  114.1958, 114.2408, 115.0983, 114.323, 112.1833, 107.9729, 95.43396,
    79.00027, 86.04683, 75.42306, 71.17786, 68.58025, 71.90591, 72.90392,
    66.97495, 56.87499, 58.1212, 58.3528, 58.30587, 60.62272, 62.62082,
    60.645, 57.02224, 53.79269, 51.86886, 46.52438, 40.556, 41.37979,
    40.59073, 39.11465,
  104.7053, 104.4786, 103.7839, 102.0637, 99.84838, 99.56402, 99.36178,
    99.49075, 91.66953, 91.9458, 96.80919, 92.78271, 90.14053, 90.13028,
    82.28601, 70.29967, 67.55861, 71.04263, 72.99384, 67.18994, 59.69049,
    54.31982, 50.42855, 44.5021, 41.38918, 41.03637, 39.95716, 39.38158,
    39.47242, 38.86335,
  79.7635, 76.23917, 78.19934, 78.5116, 79.2888, 80.67822, 83.75273,
    82.52071, 79.36427, 79.88553, 77.19704, 73.76489, 75.41331, 76.75475,
    77.24582, 75.26491, 69.6168, 66.85351, 65.17313, 60.2784, 50.33223,
    48.53745, 43.72476, 41.57694, 41.30371, 40.68352, 39.78276, 38.92474,
    38.3858, 38.01772,
  71.19562, 73.15604, 73.83216, 73.23053, 72.33936, 73.47125, 74.75356,
    71.16058, 66.55008, 63.99192, 63.79298, 61.76147, 60.31111, 63.61982,
    61.973, 61.88481, 62.35125, 58.06644, 55.37517, 50.82503, 44.50645,
    44.74853, 42.13926, 41.30562, 41.10998, 40.58506, 39.78088, 39.09356,
    38.48684, 38.0032,
  62.20988, 61.18938, 61.57125, 62.61916, 63.65055, 64.64965, 65.67221,
    66.81234, 65.82641, 63.31306, 59.68541, 63.63313, 67.86871, 64.06835,
    59.69575, 57.6761, 55.89305, 54.23789, 53.39296, 50.68269, 44.78286,
    45.02517, 42.57201, 41.28105, 40.88412, 40.75022, 39.49796, 38.40021,
    38.16203, 37.94398,
  59.53563, 60.13673, 59.1279, 60.24111, 61.37409, 62.86502, 64.01015,
    65.57057, 66.51376, 65.60542, 68.87521, 72.17476, 71.38279, 69.49947,
    64.4121, 60.11652, 56.54211, 55.87867, 56.78968, 52.70455, 45.54169,
    44.7916, 42.98387, 41.9976, 40.63468, 39.87415, 39.14342, 37.96338,
    37.8512, 37.7298,
  68.87785, 64.19284, 57.42103, 54.50401, 56.35808, 56.88366, 57.96094,
    59.16526, 59.36473, 61.26615, 64.64938, 63.84604, 59.98824, 61.532,
    61.98129, 64.55269, 69.69993, 73.31918, 71.6225, 64.0662, 53.29688,
    47.06192, 43.85379, 42.58554, 40.77771, 39.67546, 38.97997, 38.08479,
    37.80012, 37.72989,
  65.17099, 60.65159, 54.48344, 51.22994, 52.97953, 53.85608, 54.93707,
    56.08011, 57.89708, 61.23008, 61.81459, 57.48642, 57.59641, 57.08944,
    56.53069, 57.13167, 59.96703, 63.73591, 64.63242, 62.57643, 57.23321,
    50.67797, 45.79043, 44.15181, 42.57064, 40.4298, 39.25956, 38.20718,
    37.76097, 37.74265,
  60.91435, 56.95079, 50.85426, 47.87537, 48.92362, 49.56613, 50.46184,
    51.49008, 53.32961, 55.25121, 53.35827, 50.60573, 52.9877, 52.8517,
    51.81513, 51.4579, 52.32608, 53.63534, 54.66109, 53.80682, 53.10005,
    52.63216, 49.52118, 46.66876, 44.09542, 41.24632, 39.3121, 38.2956,
    37.78074, 37.7591,
  59.61432, 56.1848, 50.16445, 47.47577, 47.97741, 47.16644, 47.86721,
    48.48328, 50.59146, 51.15989, 47.76863, 46.1153, 47.82488, 48.22116,
    48.15703, 48.49129, 48.63916, 49.19648, 50.13192, 50.3786, 50.24119,
    49.95631, 50.003, 49.15344, 46.01753, 41.78886, 39.55978, 38.66585,
    37.88709, 37.74555,
  62.25733, 60.82247, 53.84897, 51.5334, 53.03764, 52.86713, 51.52665,
    49.62236, 50.02523, 48.92553, 45.71407, 46.41762, 47.40107, 48.08977,
    47.90457, 48.48444, 48.67778, 47.84436, 47.8382, 47.90028, 47.68176,
    47.05848, 46.37852, 46.957, 47.18488, 43.63897, 40.58917, 39.81997,
    38.61599, 37.83009,
  68.52641, 68.05711, 63.36311, 61.63764, 61.38012, 60.26618, 60.43719,
    59.68671, 60.96478, 58.08371, 54.76995, 56.4287, 57.72909, 58.31014,
    57.15111, 56.13177, 55.19176, 53.44334, 51.36085, 50.18148, 49.08198,
    48.06439, 47.08109, 46.71283, 47.7091, 47.72266, 44.7042, 41.28989,
    39.97684, 38.44774,
  71.92501, 67.76293, 61.81949, 59.42296, 59.49398, 58.93287, 60.02565,
    63.01588, 66.4539, 62.83796, 58.25074, 60.01595, 61.21288, 62.05634,
    61.39696, 60.64319, 59.0322, 57.54465, 55.357, 53.17166, 51.94997,
    50.57981, 48.34428, 46.82428, 47.61766, 49.20933, 48.84573, 44.47317,
    41.64546, 39.62906,
  75.00537, 71.68277, 66.44087, 62.1907, 60.60826, 59.99893, 62.9755,
    66.87462, 66.60114, 62.21091, 61.31971, 62.09, 62.9941, 62.50564,
    61.05537, 60.60951, 59.91183, 58.87625, 56.99651, 55.03814, 54.33241,
    52.98582, 49.60847, 47.56275, 47.87426, 48.56941, 49.09279, 45.59496,
    40.85438, 39.11411,
  76.0787, 71.65938, 66.82622, 63.57072, 61.92192, 60.34624, 63.41122,
    65.07436, 64.00119, 62.21555, 63.23363, 63.60294, 63.78749, 63.43492,
    62.47534, 61.76791, 61.3772, 60.76939, 59.29264, 58.15217, 58.63497,
    58.93658, 56.53611, 53.20257, 52.19527, 52.43115, 53.03224, 49.31884,
    41.52704, 38.21091,
  73.54516, 70.63414, 67.66864, 67.1411, 67.11994, 65.72288, 64.88857,
    63.30696, 60.9418, 61.51646, 62.23632, 63.21135, 64.17767, 64.62906,
    64.70755, 64.1797, 63.07454, 62.11245, 61.35004, 60.88094, 59.64378,
    57.11742, 54.01074, 52.19687, 51.67743, 52.12588, 52.01334, 52.07019,
    47.72362, 39.92328,
  60.79619, 60.561, 61.34478, 62.2295, 64.01736, 65.70123, 62.23241,
    55.62047, 53.86455, 54.5178, 54.10503, 54.47073, 55.43728, 56.34289,
    57.06858, 57.39988, 56.74845, 55.7463, 53.60868, 51.53434, 50.38846,
    49.08359, 47.57745, 46.44715, 46.5192, 46.33653, 45.66838, 44.52949,
    43.81339, 40.97245,
  54.84034, 55.23572, 55.25139, 54.87978, 56.85309, 60.85628, 60.92728,
    54.24914, 51.63893, 53.78199, 55.14204, 56.25769, 56.13468, 54.50504,
    52.42056, 51.21099, 48.39594, 46.1186, 45.8875, 44.90783, 43.77001,
    43.78883, 43.83654, 43.66366, 43.40243, 43.27098, 42.48248, 41.0439,
    39.45031, 37.95063,
  40.77556, 40.76947, 40.82731, 40.89202, 40.89886, 40.98538, 41.13519,
    41.38885, 41.7032, 42.21488, 43.11745, 42.94172, 41.52355, 41.95182,
    42.04752, 41.53148, 41.52757, 41.72038, 42.05579, 42.79494, 43.13519,
    42.44947, 42.81072, 44.2365, 45.70026, 46.19557, 48.11677, 49.26601,
    43.60261, 41.64738,
  41.73039, 41.80492, 41.46968, 41.85382, 41.69378, 41.69879, 42.00809,
    42.35411, 42.77188, 43.23712, 43.79184, 44.27851, 44.39617, 43.51598,
    42.9046, 43.0993, 42.49824, 43.01464, 43.8205, 44.49046, 44.80091,
    45.42936, 47.45612, 51.7784, 55.69687, 52.38092, 47.26339, 49.77544,
    44.31221, 42.23757,
  41.32193, 41.27877, 41.29574, 41.36715, 41.42992, 41.63314, 41.89666,
    42.23751, 42.63616, 42.98914, 43.41007, 44.05453, 44.61889, 45.41965,
    46.01978, 45.60978, 46.69631, 48.4405, 50.17716, 53.2267, 58.72482,
    65.31151, 67.34258, 65.00677, 62.78771, 58.41337, 54.07872, 49.03357,
    44.41197, 42.93177,
  42.28379, 42.78024, 43.60719, 44.48616, 45.3109, 46.20567, 46.46764,
    46.52444, 46.92944, 47.46851, 48.02438, 48.9578, 49.58132, 49.92847,
    52.45481, 54.46157, 54.6012, 55.59648, 59.45304, 64.38671, 71.17137,
    71.44637, 65.26103, 65.04859, 61.67663, 60.07179, 58.37023, 50.56285,
    43.85404, 41.89026,
  45.74935, 46.034, 47.11183, 47.86787, 48.28633, 48.30254, 48.26488,
    48.06595, 48.49674, 48.6698, 48.64381, 50.05321, 51.47256, 53.01445,
    55.20479, 57.71742, 58.58328, 58.84439, 62.46317, 67.40425, 66.92452,
    58.50867, 56.13694, 58.95815, 60.6895, 60.44771, 59.4982, 64.28874,
    62.00903, 48.29617,
  47.12746, 48.06034, 49.3934, 50.59648, 50.12495, 49.84558, 51.54779,
    52.90762, 54.94135, 58.45554, 64.02216, 74.24818, 82.93317, 80.85318,
    81.9257, 84.06082, 81.64359, 76.31984, 69.96036, 67.17951, 60.52618,
    53.63038, 57.32123, 60.25389, 63.90571, 65.43429, 67.4919, 77.19926,
    71.2967, 46.30053,
  51.46273, 54.16647, 57.17676, 60.39388, 63.31912, 68.79446, 78.31123,
    86.91851, 89.60912, 89.16732, 88.64628, 83.58008, 75.54346, 74.90187,
    74.5845, 74.24004, 73.30075, 68.09735, 62.66166, 60.90286, 57.54,
    56.74225, 59.70262, 63.14464, 64.87933, 64.60385, 69.31679, 74.89429,
    61.81959, 40.82536,
  61.69019, 66.34961, 70.54986, 75.11746, 79.09854, 86.65391, 91.02223,
    80.29741, 72.89184, 70.82302, 66.30503, 61.52943, 58.27545, 57.93293,
    58.03262, 59.32693, 60.49747, 59.38884, 57.09463, 56.91603, 56.72211,
    57.88596, 60.65446, 63.15351, 63.00838, 64.7594, 71.03589, 69.56931,
    54.13216, 40.80754,
  68.85211, 71.62863, 73.4479, 74.78305, 76.86746, 76.76363, 66.56621,
    60.86721, 60.29121, 58.8933, 57.74518, 57.6422, 59.08393, 63.44809,
    65.53804, 61.34668, 62.4627, 64.66956, 63.93148, 61.06895, 60.25006,
    63.73197, 67.84099, 67.69569, 66.09087, 71.64275, 73.25278, 62.11229,
    43.42237, 41.49213,
  71.81642, 74.29127, 71.59102, 72.08454, 73.67408, 68.55433, 55.23376,
    59.50441, 60.44059, 63.61711, 67.35011, 71.29575, 71.54372, 70.64155,
    69.2289, 71.34552, 73.18192, 73.00263, 71.40298, 70.77519, 72.00746,
    71.20211, 68.91771, 65.35793, 69.19159, 75.68277, 68.29784, 49.13022,
    40.82627, 40.72487,
  72.82175, 72.73612, 72.87917, 73.00156, 76.82668, 72.07441, 66.29371,
    71.24158, 75.45868, 75.8036, 69.5661, 61.79433, 60.77205, 61.45445,
    62.3202, 63.82337, 65.36353, 65.79688, 65.89043, 67.6498, 71.56416,
    69.26832, 62.72107, 61.54041, 66.45226, 64.68447, 50.6711, 41.01469,
    41.33509, 40.61826,
  80.45465, 74.86035, 82.14029, 87.28674, 83.96533, 75.1252, 77.33504,
    71.63094, 66.19957, 64.41051, 59.7089, 57.28394, 59.34912, 59.871,
    58.96556, 59.66281, 59.24052, 59.4154, 59.68204, 61.61195, 65.78672,
    65.08997, 60.88491, 65.69126, 66.87003, 54.92873, 41.62053, 43.16327,
    41.79975, 41.01395,
  100.73, 103.6883, 106.394, 106.4372, 104.6177, 100.8196, 83.65723,
    71.61982, 76.93099, 69.10136, 65.4566, 64.34898, 67.8618, 69.28576,
    65.31436, 57.21299, 58.4631, 58.91145, 59.43438, 62.33645, 65.59698,
    65.34171, 62.72916, 58.90142, 55.63779, 49.12119, 42.87003, 44.18198,
    43.19491, 41.878,
  104.4864, 105.66, 104.4731, 100.8283, 97.60394, 95.34517, 93.9278,
    93.21984, 85.58242, 85.97772, 90.64156, 87.19795, 84.83236, 84.36042,
    78.29308, 68.041, 66.48759, 71.51047, 74.51148, 70.80859, 65.71742,
    60.91122, 55.658, 48.84336, 45.04292, 44.18875, 43.0946, 42.56233,
    42.47941, 41.76478,
  98.62041, 94.33577, 91.24196, 87.64085, 86.50597, 89.6256, 94.78661,
    91.58697, 86.57632, 86.7739, 83.7997, 79.31404, 79.0479, 80.96706,
    80.56433, 78.90005, 75.13348, 73.05499, 71.58566, 66.35835, 56.14627,
    52.6405, 46.96978, 43.92203, 43.69477, 43.39928, 42.63876, 41.83699,
    41.38466, 40.99539,
  84.39598, 84.80779, 85.14915, 83.9353, 82.78526, 83.71927, 84.34594,
    80.40068, 75.67035, 72.45589, 71.16473, 68.57396, 68.39584, 71.29773,
    69.2035, 68.25925, 67.45149, 62.59711, 59.2353, 54.05036, 47.70631,
    47.01497, 44.15717, 43.39142, 43.47371, 43.2214, 42.52964, 41.85597,
    41.29344, 40.89834,
  74.62814, 73.30077, 72.43998, 71.73126, 71.10603, 70.38731, 70.14037,
    70.31975, 68.64042, 66.07269, 62.90276, 65.54912, 69.42403, 66.71172,
    62.11217, 59.96116, 57.86951, 55.67316, 54.55531, 51.91405, 46.70871,
    46.81978, 44.69038, 43.48646, 43.36166, 43.43028, 42.37538, 41.40597,
    41.08816, 40.85954,
  63.6983, 63.7199, 62.78471, 63.17579, 63.56725, 64.55672, 65.48354,
    66.55447, 66.56995, 65.18961, 67.57929, 70.21714, 69.34563, 66.84111,
    62.17071, 58.13228, 54.80387, 54.31139, 55.37798, 52.61964, 47.19057,
    46.78668, 45.18443, 44.22934, 43.21513, 42.60763, 41.95934, 40.97731,
    40.82047, 40.70893,
  69.68217, 66.23643, 60.19951, 57.38675, 58.75151, 58.86698, 59.50568,
    60.0023, 59.57548, 60.75346, 63.25755, 61.67837, 57.253, 57.35894,
    56.43767, 57.99796, 62.62468, 67.02124, 67.1004, 61.8889, 53.64163,
    48.85839, 46.0431, 44.8656, 43.24867, 42.36455, 41.78903, 41.0391,
    40.7624, 40.70018,
  69.07736, 64.14262, 57.50363, 53.87442, 54.86546, 54.80832, 54.99039,
    55.32558, 56.45094, 59.36227, 60.02488, 56.59702, 56.75686, 56.65853,
    56.63132, 58.10248, 61.61151, 65.45913, 65.72623, 62.89062, 57.53717,
    51.64101, 47.43156, 46.03167, 44.61427, 43.01331, 42.05896, 41.15329,
    40.76638, 40.71309,
  66.02445, 61.92366, 55.43571, 52.23766, 53.04927, 53.30202, 53.76715,
    54.6227, 56.50827, 58.7965, 57.72095, 55.84181, 58.07994, 57.99961,
    57.14233, 56.78314, 57.18669, 57.64067, 57.40425, 55.34952, 53.90771,
    53.04946, 50.42478, 47.99533, 45.86378, 43.69437, 42.08958, 41.19237,
    40.77423, 40.74735,
  64.18, 61.14173, 55.22984, 52.94663, 53.76212, 53.52077, 54.53111,
    55.39664, 57.40826, 57.98242, 55.04253, 53.47567, 54.47537, 53.94413,
    53.1129, 52.752, 52.26641, 52.11486, 52.32257, 52.12505, 51.86137,
    51.74274, 51.74914, 50.28998, 47.45176, 44.20199, 42.23925, 41.47454,
    40.81931, 40.71338,
  62.38934, 60.91082, 55.00639, 53.41457, 55.27819, 55.71489, 55.08345,
    53.83578, 54.03356, 52.73837, 49.60688, 49.66273, 50.16065, 50.23237,
    49.89468, 50.45519, 50.72926, 50.25463, 50.30501, 50.27627, 50.0081,
    49.5969, 48.9654, 48.53123, 48.1659, 45.29912, 42.84679, 42.20567,
    41.2966, 40.77061,
  64.36064, 64.08446, 59.96623, 58.5928, 58.72945, 57.576, 57.31806,
    56.64198, 57.49262, 55.13317, 52.39458, 53.85448, 55.14152, 55.74902,
    55.21917, 55.12141, 55.08967, 53.87261, 52.13019, 51.01469, 50.26098,
    49.58064, 48.48896, 47.81056, 48.46459, 48.4613, 45.90451, 43.13237,
    42.24826, 41.23783,
  67.63861, 64.70497, 59.06828, 56.74374, 56.6049, 55.80153, 56.48105,
    58.94106, 62.10242, 59.5014, 56.13963, 57.9681, 59.34324, 60.06085,
    59.59693, 59.46645, 58.76143, 57.76694, 55.8823, 54.25981, 53.35085,
    52.05006, 49.91702, 48.54692, 49.35132, 50.65566, 49.77966, 45.83032,
    43.76277, 42.25573,
  69.27293, 66.8501, 61.7029, 58.20534, 57.23929, 56.84056, 59.5408,
    63.72443, 64.45689, 60.86264, 60.0377, 61.18781, 62.38378, 62.0443,
    60.63334, 60.45709, 60.07939, 59.07629, 57.50911, 56.1306, 55.33632,
    53.7531, 50.80697, 49.29357, 49.68356, 50.12978, 50.49321, 47.36906,
    43.3799, 41.891,
  70.52733, 67.66481, 63.19936, 59.93552, 58.82893, 57.71191, 60.61687,
    62.78143, 62.30964, 60.54575, 61.23056, 61.99875, 62.61817, 62.164,
    60.88443, 60.5154, 60.44192, 59.7809, 58.47439, 57.48891, 57.54524,
    57.34203, 55.64237, 53.53186, 52.62234, 52.58157, 53.3798, 50.28434,
    43.67053, 41.0482,
  72.0476, 69.46695, 66.05537, 64.76197, 64.71558, 63.84627, 63.68802,
    62.98691, 61.11353, 61.20362, 61.78996, 62.71935, 63.77787, 63.98223,
    63.81296, 63.72913, 63.3847, 62.57532, 62.11176, 61.9086, 60.68973,
    58.36544, 55.55761, 53.81182, 53.18898, 53.23642, 53.30202, 53.01418,
    48.81602, 42.36092,
  64.71937, 64.27795, 64.46658, 64.87562, 66.46898, 68.07651, 65.53584,
    60.31813, 58.93818, 59.32228, 59.0031, 59.52896, 60.64166, 61.89394,
    62.84783, 63.20637, 62.54835, 61.24031, 59.11823, 56.99533, 55.41332,
    53.67973, 51.83585, 50.445, 50.14733, 49.90315, 49.25674, 47.82884,
    46.48447, 43.48444,
  60.82462, 61.33587, 61.55342, 61.11193, 62.85027, 66.37714, 66.25638,
    60.60213, 58.31308, 59.7453, 60.51057, 61.29632, 61.20987, 60.08429,
    58.34028, 56.9533, 54.39507, 52.00608, 51.13764, 49.7167, 48.3618,
    47.93218, 47.67569, 47.27161, 46.82565, 46.53765, 45.6722, 44.22134,
    42.70005, 41.10454,
  38.85304, 38.79264, 38.80592, 38.79992, 38.77382, 38.79248, 38.86651,
    39.02472, 39.22632, 39.53403, 40.13375, 40.14607, 39.17033, 39.40372,
    39.49669, 39.18727, 39.16968, 39.25162, 39.41981, 39.88624, 40.10038,
    39.48934, 39.49359, 40.26311, 41.32835, 41.9396, 43.25798, 44.6498,
    40.94229, 39.53569,
  39.39599, 39.41045, 39.13428, 39.34137, 39.15807, 39.11918, 39.34682,
    39.63926, 39.9926, 40.36073, 40.76221, 41.09176, 41.21506, 40.65141,
    40.02872, 40.18855, 39.73793, 39.94928, 40.25138, 40.34213, 39.81758,
    39.55562, 41.17992, 45.4066, 49.71658, 47.66045, 43.14569, 45.65337,
    41.49074, 39.99655,
  39.48144, 39.38309, 39.32734, 39.28955, 39.20904, 39.28889, 39.43676,
    39.61634, 39.76961, 39.94586, 40.19955, 40.57383, 40.87326, 41.06662,
    41.00716, 40.23798, 40.38489, 40.93951, 41.37651, 43.16989, 47.82473,
    55.01742, 59.02049, 58.53791, 57.30054, 52.85299, 49.3529, 45.23689,
    41.59071, 40.55472,
  39.518, 39.53099, 39.8296, 40.19766, 40.49347, 41.00086, 41.18754,
    41.22689, 41.55019, 42.05345, 42.42521, 42.80276, 42.75313, 42.32498,
    43.34813, 44.12312, 43.96935, 44.65516, 48.26989, 54.21445, 62.97254,
    66.13852, 60.94541, 60.29597, 56.66226, 55.40187, 54.45248, 46.84715,
    40.60526, 39.50159,
  40.58399, 40.55964, 41.43157, 42.16447, 42.70307, 43.08574, 43.29434,
    43.14561, 43.11375, 42.43472, 41.20043, 40.68674, 40.58984, 41.54132,
    43.34288, 45.88477, 48.05928, 50.73201, 56.57604, 63.44989, 64.97783,
    56.86051, 52.49, 54.39074, 55.05636, 54.84936, 54.48869, 59.31767,
    58.17893, 46.00282,
  41.95211, 42.70688, 43.62706, 44.10635, 43.07986, 41.70554, 41.16769,
    40.50077, 40.54134, 42.27953, 46.06976, 54.9047, 64.29669, 64.87114,
    68.3762, 72.24905, 72.8013, 71.71931, 68.17085, 65.27218, 57.36361,
    48.2058, 50.93995, 53.46149, 56.74158, 58.75884, 61.51246, 71.69833,
    69.02612, 45.09985,
  42.52294, 42.88119, 43.2937, 43.78753, 44.14256, 46.64905, 53.91806,
    63.63809, 68.98898, 71.58771, 75.28038, 74.57968, 70.23987, 72.14501,
    73.79652, 74.37543, 73.86079, 68.05748, 60.66259, 56.38407, 51.53339,
    50.27905, 53.96675, 57.65994, 60.49089, 61.46794, 66.13028, 71.82198,
    60.2646, 38.93888,
  43.33915, 45.23498, 48.28694, 52.74536, 58.33549, 68.85249, 78.61693,
    74.13528, 70.70851, 71.83362, 69.87376, 65.92791, 62.80677, 62.29026,
    61.18599, 60.59956, 59.28501, 55.91541, 52.40045, 51.83886, 51.89533,
    53.61335, 56.71179, 59.57591, 60.29169, 62.14007, 67.63856, 66.35789,
    51.98821, 38.83175,
  50.81558, 55.56387, 60.48366, 66.02301, 73.13774, 77.70105, 70.72915,
    65.22991, 64.58792, 62.85941, 60.59203, 58.98678, 58.84929, 60.4781,
    60.66976, 56.23054, 56.03299, 57.52562, 57.52683, 55.66243, 55.31286,
    58.54537, 62.45465, 62.99169, 61.93893, 67.81299, 70.67419, 60.5521,
    41.41045, 39.3551,
  63.036, 69.62962, 70.13988, 73.61227, 77.0119, 72.70428, 57.21273, 59.2667,
    58.76339, 60.1772, 62.55373, 65.11761, 64.50519, 63.05509, 61.22092,
    62.02766, 63.78118, 64.50571, 63.96624, 63.72659, 65.05647, 65.07031,
    64.06502, 61.10338, 64.64313, 72.21391, 67.35811, 47.87262, 38.93114,
    38.8861,
  71.67694, 75.00802, 74.13167, 72.23897, 73.33825, 65.77428, 58.17547,
    63.65498, 67.6774, 69.47655, 65.38045, 58.68312, 57.26525, 57.17908,
    57.39693, 58.98948, 60.47098, 61.09548, 61.73167, 63.64426, 67.32437,
    65.66312, 60.57614, 60.21896, 65.75198, 64.86823, 50.51332, 39.17895,
    39.38828, 38.7061,
  76.01884, 67.38833, 69.90041, 73.10344, 71.72817, 66.25976, 72.30708,
    68.99325, 63.36843, 62.90065, 57.562, 54.25976, 56.16871, 56.73067,
    55.87322, 57.21393, 57.29658, 57.67804, 58.03426, 59.67222, 63.3217,
    62.86097, 59.71645, 64.45417, 66.03853, 54.50896, 39.67526, 40.88515,
    39.81903, 38.99491,
  87.8207, 90.08907, 94.20261, 96.73393, 97.49393, 95.7174, 80.51591,
    65.53993, 70.37678, 63.17569, 59.48962, 59.76109, 64.2728, 66.30383,
    63.16902, 55.22939, 56.26288, 56.58188, 56.90253, 59.33746, 63.08389,
    64.33371, 63.2612, 59.52203, 54.59446, 47.08888, 40.27432, 42.08166,
    40.86877, 39.7981,
  94.33159, 99.17087, 101.0069, 98.92609, 95.6845, 91.5877, 86.07607,
    84.88052, 76.90851, 77.05894, 82.81, 81.60288, 80.54036, 80.62622,
    74.25227, 63.22177, 61.89476, 67.32765, 71.18515, 68.85313, 65.76197,
    61.6598, 55.52222, 48.24507, 43.5069, 42.00208, 40.99765, 40.69902,
    40.3716, 39.75077,
  97.58976, 98.18363, 94.95123, 88.81683, 82.20999, 82.6621, 88.62747,
    87.76009, 82.94019, 83.88525, 81.57121, 76.40607, 75.87708, 77.77988,
    77.83386, 77.65077, 74.68428, 73.94977, 72.39742, 67.22579, 56.96827,
    52.35917, 45.59671, 41.73705, 41.54514, 41.31849, 40.65227, 39.89315,
    39.48776, 39.10393,
  92.04331, 87.14703, 83.42973, 80.48244, 79.95598, 82.88968, 84.88274,
    81.30023, 76.7841, 72.56606, 70.11825, 67.9708, 68.85767, 73.13564,
    72.42881, 71.47169, 70.66115, 65.29849, 60.12819, 53.53725, 46.85093,
    45.01858, 41.7544, 41.0207, 41.33021, 41.10833, 40.41278, 39.78736,
    39.30684, 38.97789,
  80.1725, 77.15662, 76.76933, 76.73209, 76.23476, 74.55105, 72.82776,
    71.75684, 69.17343, 66.3697, 64.09396, 66.6809, 70.86527, 69.70208,
    65.05035, 61.98949, 58.68557, 54.88297, 51.79783, 48.67938, 44.11689,
    43.94755, 41.98789, 41.09665, 41.00842, 41.04485, 40.24586, 39.46879,
    39.12176, 38.92929,
  71.73535, 71.91405, 70.90334, 70.06412, 68.56499, 67.57883, 67.19493,
    67.7513, 67.90817, 66.811, 68.73009, 71.2795, 70.48386, 67.10822,
    61.47749, 56.83184, 52.33931, 50.14486, 49.87268, 47.77555, 43.72248,
    43.78268, 42.32787, 41.55693, 40.95607, 40.5163, 39.94365, 39.10342,
    38.92337, 38.80661,
  77.23503, 73.87164, 67.37703, 63.42227, 64.02869, 63.93876, 64.59014,
    65.32874, 65.09727, 65.67421, 66.84925, 64.44939, 58.68398, 56.08206,
    52.81225, 52.08199, 54.42997, 57.57565, 58.29414, 55.31388, 49.69658,
    45.87909, 43.22403, 42.41817, 41.06865, 40.38055, 39.86384, 39.11397,
    38.8448, 38.7896,
  76.5537, 70.79161, 63.98917, 60.41988, 61.56791, 61.60139, 61.57699,
    61.17508, 60.94122, 61.5811, 60.11711, 54.99467, 52.63139, 50.89694,
    49.95186, 51.21973, 54.98106, 59.52551, 60.61389, 58.4636, 53.77023,
    48.32078, 44.4518, 43.41973, 42.09938, 40.89267, 40.13328, 39.24728,
    38.82173, 38.78839,
  72.27643, 67.86013, 61.47678, 58.00322, 58.40842, 57.74451, 56.98865,
    56.13346, 55.8972, 55.98233, 53.73808, 51.17774, 52.84071, 53.24149,
    53.55887, 54.54488, 55.94148, 56.59887, 55.68959, 52.76346, 50.29844,
    48.83006, 46.62797, 44.98295, 43.21948, 41.48682, 40.17882, 39.30485,
    38.83392, 38.79334,
  68.87777, 65.39857, 58.88106, 55.43044, 55.21299, 53.86464, 53.63618,
    53.45438, 54.47483, 54.95127, 53.06941, 52.5793, 54.60192, 54.9948,
    54.62156, 54.14114, 52.87441, 51.34119, 50.18863, 48.99966, 48.34643,
    48.06888, 47.99843, 46.67469, 44.43573, 41.84593, 40.36299, 39.56865,
    38.90907, 38.82455,
  65.76065, 62.98114, 56.20317, 53.577, 54.69541, 54.68282, 54.26942,
    53.73265, 54.7369, 54.52426, 52.40891, 52.8461, 53.19724, 52.64455,
    51.22449, 50.26511, 49.21417, 47.97577, 47.56731, 47.33168, 47.21334,
    46.84509, 46.11457, 45.30323, 44.85122, 42.52042, 40.54019, 40.11187,
    39.29231, 38.85205,
  65.365, 64.42364, 59.86331, 58.24274, 58.58474, 57.65582, 57.58705,
    57.4845, 59.06775, 57.53539, 54.77722, 55.34121, 55.50067, 54.70624,
    53.07574, 52.05529, 51.50838, 50.38406, 48.93964, 48.01568, 47.38943,
    46.74327, 45.51299, 44.74441, 45.02034, 44.51426, 42.55084, 40.71602,
    40.09365, 39.30796,
  68.97602, 66.44424, 60.69529, 58.0499, 57.67786, 56.80308, 57.47925,
    59.5858, 62.61541, 60.14058, 56.44523, 57.11896, 57.48492, 57.5152,
    56.50543, 55.91377, 55.01327, 53.97426, 52.04829, 50.39616, 49.55982,
    48.62111, 46.60844, 45.32403, 45.74068, 46.10611, 45.27397, 42.75693,
    41.40702, 40.2084,
  69.89093, 67.50196, 61.82168, 58.05484, 57.23279, 56.61707, 58.91309,
    62.57961, 63.42887, 59.87088, 58.73154, 59.26332, 59.96619, 59.69575,
    58.12052, 57.51718, 56.80761, 55.69458, 54.03275, 52.69236, 51.87362,
    50.26519, 47.65675, 46.35154, 46.64593, 46.30937, 46.09841, 44.11541,
    41.24742, 39.95385,
  69.48116, 66.81562, 61.97226, 58.56887, 57.97181, 57.10546, 59.61333,
    61.70154, 61.60329, 59.77217, 60.15284, 60.52811, 60.79251, 60.11009,
    58.56315, 57.57988, 57.0789, 56.19537, 55.06262, 54.17265, 53.54102,
    52.93319, 51.2879, 49.72308, 49.08737, 48.34273, 48.54715, 46.35847,
    41.25271, 39.22001,
  69.14014, 66.29942, 62.81264, 61.44809, 62.26785, 61.92717, 62.27152,
    62.16437, 60.86929, 60.64785, 60.96375, 61.18671, 61.49575, 61.33512,
    60.47765, 59.58882, 58.92762, 58.10103, 57.61774, 57.44223, 56.16989,
    54.26136, 51.98103, 50.5727, 49.9489, 49.3992, 48.86834, 48.22808,
    45.09625, 40.1482,
  62.53905, 62.11598, 62.33773, 62.9627, 64.75639, 66.41147, 64.49097,
    60.36518, 58.88602, 58.81223, 58.15865, 58.23003, 58.82462, 59.61697,
    60.16907, 60.29015, 59.65608, 58.4165, 56.5048, 54.60977, 53.07223,
    51.62922, 49.91692, 48.55847, 48.09815, 47.60139, 46.88259, 45.49588,
    43.96137, 41.23122,
  59.15631, 59.81173, 60.38036, 60.39587, 61.84422, 64.91122, 64.87699,
    59.79359, 57.58879, 58.2766, 58.69028, 59.45251, 59.50738, 58.78311,
    57.61679, 56.53371, 54.10522, 51.6587, 50.29317, 48.64897, 47.2814,
    46.77512, 46.36571, 45.77757, 45.14454, 44.61531, 43.64528, 42.25145,
    40.862, 39.33648 ;

 no2_conc_recp_ens =
  39.24281, 16.32957, 39.11094, 21.15891, 15.71463, 8.199514, 30.48344,
    83.22491, 22.54597,
  85.94411, 52.97182, 86.70657, 74.09569, 61.01787, 36.84403, 82.19931,
    80.52858, 84.78162,
  80.24696, 81.96887, 82.43535, 81.53499, 82.1398, 80.45194, 81.67593,
    75.23991, 84.88847,
  79.97185, 77.58305, 82.16718, 78.95976, 76.07831, 78.48167, 80.07261,
    86.76813, 78.92854,
  84.58956, 85.64126, 83.9413, 84.77237, 84.00996, 77.40044, 89.17546,
    78.05194, 78.45639,
  81.14112, 81.84781, 77.18153, 79.89639, 78.55714, 79.36035, 85.68592,
    73.70714, 70.50311,
  84.91205, 84.4688, 77.56792, 79.49628, 76.76386, 69.56031, 92.66521,
    91.41611, 68.62247,
  85.82564, 91.27137, 87.25397, 94.55315, 95.19691, 92.88631, 92.26633,
    74.85469, 83.19339,
  66.85131, 79.439, 63.06388, 78.14297, 64.90945, 81.52176, 67.61392,
    61.77457, 57.43208,
  46.13483, 75.10043, 44.70932, 65.30826, 54.08834, 68.06772, 48.78827,
    43.59865, 38.47776,
  43.51596, 56.43639, 42.06651, 52.33688, 37.96053, 46.94086, 45.15809,
    41.08328, 36.6632,
  32.26695, 54.89642, 31.14607, 44.0903, 29.00041, 43.41335, 34.00225,
    30.31999, 27.02503,
  23.98508, 42.85028, 22.90813, 37.36971, 17.36178, 31.842, 25.77868,
    21.88128, 19.27694,
  23.19687, 39.39555, 22.20031, 32.83269, 16.33221, 23.36798, 24.94221,
    21.49671, 18.97051,
  21.61873, 40.35111, 20.63963, 31.88234, 13.70429, 22.68604, 23.51292,
    19.32618, 16.94436,
  24.12633, 51.31326, 23.02726, 31.44651, 15.54922, 21.87194, 25.49776,
    21.59987, 18.33103,
  33.08513, 77.07889, 31.42389, 52.44142, 21.94903, 30.00189, 32.5769,
    28.68619, 22.91505,
  54.96345, 68.74166, 54.95354, 64.69698, 30.55972, 62.1544, 56.97, 46.57679,
    43.81206,
  112.848, 108.5345, 104.6554, 113.275, 62.10917, 89.61442, 116.9952,
    97.32076, 75.62785,
  99.0571, 116.3711, 88.07736, 94.38913, 94.33463, 94.08183, 110.5087,
    79.24623, 71.86822,
  85.31783, 82.88587, 76.22715, 76.81447, 73.54735, 77.01698, 90.39528,
    72.18604, 61.80579,
  84.52692, 83.83124, 70.59045, 73.20323, 72.34506, 72.87865, 82.29778,
    72.12602, 65.66008,
  86.93616, 91.63814, 71.26807, 77.09091, 67.09833, 73.70415, 78.0895,
    77.28922, 69.10799,
  84.38725, 91.06755, 68.8924, 79.47382, 66.17534, 84.79895, 75.13015,
    71.57928, 62.87773,
  30.68661, 12.3297, 30.65993, 16.22139, 11.7583, 7.36852, 23.75889,
    65.85847, 19.34895,
  69.16385, 42.09262, 69.7607, 59.03803, 48.51561, 31.32685, 65.91117,
    66.97442, 68.20583,
  67.10535, 67.15643, 69.01626, 67.55417, 67.40298, 67.99944, 68.38759,
    63.91377, 71.14106,
  66.37143, 65.53378, 68.11962, 66.37861, 64.09534, 66.09702, 67.74307,
    59.53516, 62.92219,
  65.71268, 58.15979, 57.90757, 56.81569, 55.8168, 56.05637, 64.66249,
    59.63054, 51.4019,
  62.9848, 64.40562, 63.01848, 63.05059, 62.73597, 59.69666, 66.92204,
    64.03065, 59.93224,
  66.31997, 65.99051, 66.41167, 66.95931, 66.41016, 64.18166, 70.08617,
    70.1287, 66.17212,
  70.26433, 69.99442, 69.40481, 73.30861, 72.64357, 71.74343, 71.09115,
    71.49511, 69.6329,
  62.5944, 72.09515, 60.56271, 71.56982, 65.34479, 71.47207, 68.50774,
    56.25922, 56.05387,
  48.41467, 67.37171, 47.72607, 64.19907, 49.66703, 64.8916, 51.70639,
    45.61197, 41.01498,
  35.21612, 55.56146, 35.06925, 53.15281, 38.17031, 48.93563, 38.32623,
    33.12987, 29.63481,
  27.13691, 44.22936, 26.35744, 40.25724, 25.21054, 35.93325, 29.25144,
    25.09259, 22.17528,
  21.09458, 38.86863, 20.31205, 33.11867, 15.58787, 26.79174, 23.29769,
    19.13187, 16.90736,
  18.34233, 38.14358, 17.51379, 28.37519, 11.78172, 20.96363, 20.26977,
    16.29876, 14.24788,
  18.05725, 37.73629, 17.15838, 27.41834, 10.71506, 18.0269, 19.85849,
    15.70785, 13.48912,
  19.06485, 50.13079, 17.8667, 27.904, 10.90773, 18.29242, 20.50368,
    16.59319, 13.56785,
  27.73787, 75.02687, 25.74384, 44.84813, 17.19537, 25.9696, 27.20483,
    23.64584, 17.56274,
  44.57879, 72.8909, 45.95377, 62.58308, 23.76096, 64.50678, 50.64357,
    36.22237, 37.30082,
  101.3673, 98.8565, 101.6061, 103.3783, 47.8546, 87.42657, 106.3739,
    88.32539, 70.1077,
  87.89755, 103.9559, 72.80952, 79.33427, 80.50265, 87.3148, 99.56738,
    75.01892, 53.6932,
  73.67525, 74.38046, 66.57902, 68.71878, 65.00998, 64.43863, 82.14104,
    63.41798, 50.92882,
  77.63546, 69.8847, 62.74153, 63.11673, 60.83983, 62.1026, 75.14579,
    68.40044, 55.31012,
  79.46599, 85.06323, 62.63857, 68.0958, 64.18956, 64.23256, 70.72046,
    69.58135, 59.99785,
  81.92183, 83.97999, 61.58734, 73.31532, 58.68199, 76.70007, 67.9564,
    68.21496, 57.29087,
  35.59893, 16.91916, 35.51986, 21.10933, 16.78028, 7.388491, 28.94599,
    70.68681, 19.23276,
  72.95064, 47.33387, 73.87105, 63.83132, 53.52596, 31.06109, 70.55196,
    67.72269, 71.68953,
  68.92324, 69.33916, 70.9434, 69.00872, 69.0192, 68.00694, 69.79097,
    67.18539, 70.87428,
  67.9355, 63.69492, 66.24303, 63.92025, 70.05701, 62.54668, 64.71779,
    60.65815, 58.44593,
  56.94061, 61.88028, 58.1776, 60.00415, 58.95195, 56.2938, 61.52098,
    52.25321, 55.38345,
  53.6931, 55.1888, 54.09341, 54.53763, 54.49068, 57.06235, 58.25106,
    53.8772, 53.18867,
  67.81137, 59.2364, 59.90344, 63.10411, 61.01493, 54.39633, 73.87, 74.13739,
    52.76492,
  76.02912, 76.34391, 69.33096, 80.63734, 79.66918, 77.34141, 78.23009,
    61.92971, 63.67146,
  54.79171, 76.64614, 50.90741, 69.26399, 49.14161, 72.02161, 54.68183,
    49.13536, 42.82818,
  44.4694, 61.78106, 43.2104, 57.29839, 42.5524, 55.8381, 46.8408, 41.13483,
    36.57704,
  33.96842, 52.26071, 33.13189, 48.2948, 32.99449, 45.52362, 36.13877,
    31.55415, 28.40153,
  26.38601, 43.67479, 24.92654, 38.0889, 21.69327, 35.11806, 27.675,
    24.13936, 21.49503,
  19.57631, 33.8445, 18.23234, 31.76168, 12.49699, 25.21275, 21.14187,
    16.98482, 15.29809,
  22.29103, 35.62217, 21.2145, 28.94216, 15.06716, 18.85502, 23.60435,
    19.77128, 17.88773,
  22.68794, 39.90739, 21.86782, 30.44005, 15.16587, 21.51112, 24.52099,
    20.20962, 18.27827,
  27.46235, 53.85854, 26.21493, 33.35944, 19.14556, 23.778, 27.97837,
    24.82302, 20.80276,
  32.56239, 79.19848, 31.05387, 51.28608, 21.9783, 32.75383, 33.50197,
    28.6367, 23.95336,
  45.30147, 71.72462, 46.985, 62.93553, 25.49008, 65.29132, 53.24737,
    36.71515, 42.59597,
  107.9546, 99.63386, 103.7313, 108.0642, 43.34944, 89.21758, 115.9645,
    90.86785, 74.10474,
  98.81201, 117.7983, 77.86977, 96.33399, 69.91386, 94.57892, 98.0898,
    84.92195, 71.16356,
  80.43217, 92.35472, 67.30342, 72.26904, 75.81868, 73.71729, 84.40873,
    68.7505, 60.38478,
  79.25672, 87.61423, 61.31729, 69.36868, 65.30374, 67.10172, 72.97699,
    68.6452, 58.69723,
  80.22624, 83.44161, 63.14824, 73.01849, 55.40489, 75.63802, 69.51896,
    69.93386, 55.003,
  74.93463, 80.07128, 66.67047, 74.30121, 58.17641, 80.92261, 72.26804,
    66.5578, 53.23326,
  26.95305, 7.119063, 27.0634, 11.37988, 6.745733, 6.130392, 19.63688,
    64.7092, 15.8778,
  66.56714, 38.86345, 67.48846, 57.03397, 45.65199, 27.89702, 63.53453,
    57.95906, 65.91235,
  56.23025, 61.02663, 58.54482, 59.05829, 60.42937, 62.68132, 58.45456,
    51.73155, 61.81127,
  51.92426, 54.32479, 54.2306, 53.71386, 52.5548, 57.9109, 54.05716,
    50.94233, 54.56479,
  52.39023, 52.32361, 53.7527, 52.81704, 50.85582, 52.77263, 55.43585,
    53.52678, 53.19908,
  60.43183, 56.97443, 60.37873, 58.7583, 55.47502, 55.04525, 63.30087,
    65.09292, 58.7295,
  61.87544, 66.12523, 62.2458, 63.69972, 65.74121, 64.70272, 68.58321,
    64.41948, 63.30456,
  65.03912, 64.81232, 64.18105, 68.71154, 66.93838, 67.20782, 66.24061,
    69.91595, 64.73177,
  51.75903, 69.49172, 50.9664, 69.60679, 61.48865, 68.31284, 62.08033,
    44.73823, 50.16441,
  40.01011, 59.04537, 38.9316, 53.18284, 38.0373, 53.97196, 42.75164,
    37.47793, 32.38092,
  34.34415, 49.13212, 33.75363, 47.45271, 31.71303, 41.40653, 37.33067,
    32.32955, 28.32812,
  25.51551, 46.92263, 24.54278, 38.36422, 23.25251, 35.55849, 27.65954,
    23.91032, 20.7785,
  21.48863, 38.62211, 20.30159, 33.49557, 15.30061, 26.01786, 23.36147,
    19.54073, 17.09434,
  20.25713, 37.26475, 18.89875, 31.01234, 13.35779, 21.18606, 21.75427,
    18.21848, 16.02712,
  20.10013, 38.32019, 18.5239, 30.06491, 12.09454, 19.98916, 21.70603,
    17.63089, 15.37334,
  23.2226, 51.14721, 21.3513, 31.24689, 14.74251, 20.18779, 23.53905,
    20.47442, 16.46956,
  28.01364, 76.45933, 25.47098, 44.3571, 16.04572, 27.74525, 28.70011,
    22.55277, 18.92451,
  42.25581, 65.3409, 42.33096, 60.93998, 21.97726, 55.96358, 47.08779,
    34.08526, 34.22657,
  114.0894, 98.7503, 102.5443, 110.5769, 44.02725, 80.94949, 121.3382,
    91.25765, 68.9482,
  97.51505, 120.6503, 80.37849, 91.30595, 80.30768, 88.36859, 104.0674,
    83.05035, 66.14744,
  82.59921, 84.9929, 71.91276, 74.0973, 71.52849, 72.92699, 87.83609,
    72.9631, 58.82943,
  84.13082, 87.72395, 69.74864, 73.65452, 71.2664, 69.52666, 79.41427,
    76.14223, 65.57655,
  81.96664, 93.9247, 65.09779, 77.79596, 63.18715, 81.64801, 73.9799,
    69.62388, 61.03637,
  76.67582, 83.55087, 63.6137, 72.12672, 57.37471, 81.00591, 70.03235,
    65.74014, 52.21938,
  31.94525, 17.09539, 32.10018, 20.59247, 16.72886, 6.994177, 27.02182,
    59.50711, 17.70185,
  63.64368, 40.73048, 64.09897, 54.45755, 46.12275, 27.5674, 60.01668,
    65.66547, 61.8409,
  70.5938, 64.49068, 71.5931, 67.15936, 65.91481, 61.53503, 69.25407,
    68.31409, 70.76602,
  70.44604, 62.14497, 63.90114, 62.03183, 71.57158, 61.81033, 60.10682,
    53.69668, 57.69718,
  61.57814, 52.69732, 51.8917, 51.53976, 50.93441, 49.21074, 55.6847,
    48.28053, 45.39714,
  68.25157, 60.93741, 58.1972, 56.66193, 50.07636, 46.98098, 70.16285,
    65.04034, 46.04281,
  72.7756, 73.21976, 65.48464, 66.81348, 63.33824, 57.76333, 82.39737,
    77.19621, 57.34759,
  78.21124, 80.97961, 75.91147, 84.28589, 84.72513, 81.99832, 81.96545,
    65.06284, 72.12334,
  55.28559, 76.31508, 51.74846, 72.2738, 53.32347, 76.98265, 57.57408,
    49.83456, 46.47223,
  43.15131, 64.6414, 41.96008, 57.32415, 42.76118, 58.10044, 46.36324,
    40.45025, 35.6466,
  36.7737, 53.34032, 36.1525, 48.95958, 34.13894, 45.20789, 39.50606,
    34.48668, 30.77255,
  27.94857, 50.69483, 26.69427, 41.65869, 24.53725, 39.0098, 29.83963,
    25.62629, 22.83347,
  23.10378, 41.08727, 21.78185, 34.0914, 16.21981, 28.1892, 25.08889,
    20.53892, 18.60502,
  19.77773, 40.87145, 18.48143, 30.91504, 12.36001, 22.24038, 21.97109,
    17.4147, 15.97397,
  22.5309, 40.58069, 20.84167, 29.88156, 14.20201, 19.36367, 22.93135,
    19.60016, 16.33195,
  26.3996, 48.41107, 23.56579, 33.39552, 17.20345, 21.65441, 25.18443,
    22.97266, 17.94151,
  33.08838, 82.42433, 29.18054, 41.9957, 22.11672, 30.56922, 30.92027,
    28.66768, 21.35453,
  55.40355, 76.49535, 53.63919, 72.49756, 27.85151, 59.07769, 58.70369,
    44.8499, 43.85159,
  134.9683, 119.813, 113.271, 123.5499, 60.67982, 90.81255, 140.8276,
    100.2884, 80.38766,
  100.2488, 121.3082, 86.17896, 89.51692, 92.23961, 95.88968, 112.3575,
    82.09541, 68.2775,
  81.67938, 83.66985, 74.00305, 75.57057, 72.36673, 77.01357, 90.36626,
    67.99011, 57.93584,
  75.15325, 74.58586, 62.58765, 64.34844, 64.07585, 67.2812, 77.13043,
    63.24133, 54.10165,
  76.12827, 81.98558, 58.66087, 63.96632, 60.38304, 61.72338, 66.47717,
    66.89291, 56.45501,
  74.52663, 84.85918, 56.16141, 68.70158, 53.07862, 75.27498, 61.58125,
    61.06512, 50.84466,
  26.91366, 11.96891, 27.30734, 15.21408, 11.48351, 8.046144, 21.6785,
    54.64438, 18.2498,
  58.06599, 36.22455, 58.76443, 49.7264, 42.00073, 28.34892, 54.92392,
    56.29293, 57.58769,
  59.49495, 56.956, 61.29993, 58.06349, 57.67128, 58.37322, 59.09648,
    61.39186, 61.40951,
  61.48941, 61.80869, 63.5906, 62.7953, 61.2111, 60.31546, 63.86954,
    59.32549, 60.71309,
  68.84653, 61.50679, 66.43208, 64.99072, 61.06197, 58.52757, 68.54863,
    70.49769, 59.64539,
  73.89382, 77.2316, 73.94267, 75.01888, 71.4047, 67.69566, 80.05711,
    71.82122, 67.44164,
  66.92695, 71.66125, 67.25406, 68.94653, 71.61772, 69.66998, 71.63348,
    69.54279, 66.74518,
  67.39283, 70.44828, 67.7232, 72.57243, 73.68369, 72.22783, 70.31628,
    64.58032, 69.02787,
  58.34627, 66.66293, 53.69485, 65.65344, 57.80481, 66.83799, 57.2936,
    53.51839, 49.32643,
  48.44401, 66.64011, 46.20802, 58.29402, 47.02502, 58.89295, 49.29162,
    46.1053, 40.61309,
  38.50586, 55.44648, 37.5686, 51.17445, 38.88898, 48.41356, 40.32547,
    36.89069, 31.94628,
  34.0068, 49.45416, 32.65685, 43.50868, 29.71511, 38.95076, 35.40322,
    32.23335, 28.33348,
  27.83788, 43.61306, 26.95741, 39.33125, 21.87826, 33.59519, 29.77141,
    26.08469, 23.17332,
  25.20235, 44.01621, 24.01262, 35.25653, 17.94704, 27.85907, 26.38534,
    22.82608, 20.45884,
  24.47064, 43.27288, 23.27618, 34.63822, 16.58744, 24.76477, 25.99047,
    21.9612, 19.5169,
  29.04637, 59.49047, 27.80066, 36.49979, 20.47348, 26.83485, 30.17118,
    26.28072, 23.08061,
  33.72969, 82.64853, 31.72226, 57.67258, 22.2368, 36.27443, 34.97055,
    28.89464, 25.14038,
  52.92536, 76.69916, 51.66935, 64.42883, 31.73703, 72.80794, 56.43991,
    44.94683, 43.2917,
  117.3748, 110.306, 105.3435, 120.265, 54.97116, 91.43961, 127.4676,
    93.09413, 75.62931,
  99.14135, 126.7563, 82.14453, 92.63179, 88.74275, 99.83951, 106.699,
    85.42265, 68.5796,
  83.65082, 89.13232, 72.19487, 77.33143, 75.71352, 77.63158, 90.83968,
    69.05687, 62.42908,
  81.7578, 85.86821, 64.6888, 69.31566, 68.51413, 67.45598, 76.01761,
    69.27982, 61.79669,
  83.729, 91.4055, 66.88164, 75.56612, 59.76129, 77.32034, 74.20594,
    72.14912, 61.83104,
  89.43034, 89.29721, 73.43446, 80.60945, 65.46944, 84.92871, 77.3056,
    77.93029, 61.98852,
  31.69377, 16.6439, 32.1439, 20.06941, 16.38756, 7.884311, 26.5384,
    59.42526, 18.36129,
  62.78831, 40.86625, 63.76461, 54.50978, 46.50164, 28.74907, 59.7423,
    62.5732, 61.9731,
  67.19959, 62.34986, 68.76141, 64.27351, 63.19919, 62.10343, 65.85366,
    72.65906, 68.16293,
  73.16323, 67.60986, 72.51889, 70.17691, 71.96526, 63.79626, 70.1173,
    68.54007, 64.29755,
  63.9099, 66.21019, 63.21273, 64.2866, 62.86234, 60.85345, 69.99895,
    56.48174, 58.18856,
  61.95675, 60.8377, 62.10638, 61.35269, 59.92874, 60.42159, 65.58327,
    64.01528, 54.93042,
  61.18807, 65.22493, 61.55294, 62.97012, 64.37838, 59.09032, 65.59818,
    63.19045, 59.37946,
  66.2822, 64.51817, 64.41073, 67.48518, 67.3202, 66.28667, 65.29224,
    65.99203, 64.07759,
  57.40081, 71.80902, 54.4122, 71.75636, 55.67168, 70.34279, 60.0709,
    51.60734, 48.85149,
  44.42122, 65.87791, 43.11885, 60.01135, 44.72021, 59.60165, 47.48492,
    41.29211, 36.53218,
  36.20512, 52.27504, 35.54029, 50.6543, 34.51604, 45.2494, 38.89534,
    33.78772, 29.93125,
  28.34189, 45.69044, 27.11563, 40.73745, 24.24651, 37.01578, 30.10484,
    25.96439, 23.18151,
  24.15427, 36.53428, 22.88736, 35.54005, 17.16795, 27.37795, 25.98696,
    21.7479, 19.71612,
  22.85874, 40.09867, 21.46009, 33.62799, 15.64986, 23.30384, 24.78281,
    20.51551, 18.65703,
  22.71664, 40.77842, 21.41953, 31.79147, 14.98545, 21.68277, 24.69601,
    20.52308, 18.14012,
  24.77123, 53.56347, 23.31824, 32.93748, 16.36906, 22.36574, 25.94462,
    22.06595, 18.59382,
  33.71286, 80.39795, 31.3416, 49.9242, 23.23097, 31.1486, 32.86319,
    29.93114, 22.3368,
  47.95771, 75.6863, 50.04906, 70.32121, 25.29627, 66.5173, 57.11664,
    36.09285, 44.3901,
  105.0183, 104.4725, 105.0566, 106.1152, 48.45074, 89.81766, 109.5811,
    86.0322, 71.93568,
  92.38502, 112.5989, 74.44116, 85.3709, 78.93533, 90.36945, 99.47745,
    77.19547, 64.07841,
  75.15092, 79.45612, 64.06094, 66.86537, 65.86073, 68.70409, 81.27657,
    63.17996, 54.85311,
  75.26491, 79.2888, 59.69575, 63.99192, 62.13012, 62.20988, 71.38279,
    65.74888, 57.59641,
  78.90005, 86.50597, 62.11217, 72.45589, 55.23376, 74.62814, 69.34563,
    68.91771, 56.75686,
  77.65077, 82.20999, 65.05035, 72.56606, 57.21273, 80.1725, 70.48386,
    64.06502, 52.63139 ;

 dimcrs = 1 ;

 crs = "" ;

 lat =
  51.7861098779549, 51.7861349033833, 51.7861581413062, 51.7861795917181,
    51.7861992546137, 51.7862171299884, 51.7862332178379, 51.7862475181583,
    51.7862600309461, 51.7862707561984, 51.7862796939126, 51.7862868440865,
    51.7862922067185, 51.7862957818071, 51.7862975693517, 51.7862975693517,
    51.7862957818071, 51.7862922067185, 51.7862868440865, 51.7862796939126,
    51.7862707561984, 51.7862600309461, 51.7862475181583, 51.7862332178379,
    51.7862171299884, 51.7861992546137, 51.7861795917181, 51.7861581413062,
    51.7861349033833, 51.7861098779549,
  51.7951010977434, 51.795126131202, 51.7951493765815, 51.7951708338765,
    51.7951905030816, 51.7952083841922, 51.795224477204, 51.7952387821131,
    51.7952512989161, 51.7952620276099, 51.7952709681921, 51.7952781206604,
    51.7952834850131, 51.795287061249, 51.7952888493672, 51.7952888493672,
    51.795287061249, 51.7952834850131, 51.7952781206604, 51.7952709681921,
    51.7952620276099, 51.7952512989161, 51.7952387821131, 51.795224477204,
    51.7952083841922, 51.7951905030816, 51.7951708338765, 51.7951493765815,
    51.795126131202, 51.7951010977434,
  51.8040923036791, 51.8041173451711, 51.8041405980102, 51.8041620621909,
    51.804181737708, 51.8041996245568, 51.804215722733, 51.8042300322327,
    51.8042425530524, 51.8042532851892, 51.8042622286405, 51.8042693834041,
    51.8042747494783, 51.8042783268618, 51.8042801155537, 51.8042801155537,
    51.8042783268618, 51.8042747494783, 51.8042693834041, 51.8042622286405,
    51.8042532851892, 51.8042425530524, 51.8042300322327, 51.804215722733,
    51.8041996245568, 51.804181737708, 51.8041620621909, 51.8041405980102,
    51.8041173451711, 51.8040923036791,
  51.8130834957631, 51.8131085452917, 51.8131318055934, 51.8131532766626,
    51.8131729584942, 51.8131908510834, 51.813206954426, 51.8132212685181,
    51.8132337933561, 51.8132445289372, 51.8132534752587, 51.8132606323185,
    51.8132660001149, 51.8132695786465, 51.8132713679125, 51.8132713679125,
    51.8132695786465, 51.8132660001149, 51.8132606323185, 51.8132534752587,
    51.8132445289372, 51.8132337933561, 51.8132212685181, 51.813206954426,
    51.8131908510834, 51.8131729584942, 51.8131532766626, 51.8131318055934,
    51.8131085452917, 51.8130834957631,
  51.8220746739965, 51.8220997315648, 51.822122999332, 51.8221444772925,
    51.8221641654411, 51.8221820637731, 51.8221981722841, 51.8222124909704,
    51.8222250198284, 51.8222357588551, 51.822244708048, 51.8222518674049,
    51.8222572369241, 51.8222608166043, 51.8222626064446, 51.8222626064446,
    51.8222608166043, 51.8222572369241, 51.8222518674049, 51.822244708048,
    51.8222357588551, 51.8222250198284, 51.8222124909704, 51.8221981722841,
    51.8221820637731, 51.8221641654411, 51.8221444772925, 51.822122999332,
    51.8220997315648, 51.8220746739965,
  51.8310658383803, 51.8310909039916, 51.8311141792273, 51.8311356640817,
    51.8311553585498, 51.8311732626268, 51.8311893763084, 51.8312036995906,
    51.8312162324702, 51.8312269749439, 51.8312359270093, 51.8312430886642,
    51.831248459907, 51.8312520407361, 51.8312538311509, 51.8312538311509,
    51.8312520407361, 51.831248459907, 51.8312430886642, 51.8312359270093,
    51.8312269749439, 51.8312162324702, 51.8312036995906, 51.8311893763084,
    51.8311732626268, 51.8311553585498, 51.8311356640817, 51.8311141792273,
    51.8310909039916, 51.8310658383803,
  51.8400569889156, 51.840082062573, 51.8401053452801, 51.8401268370313,
    51.8401465378214, 51.8401644476457, 51.8401805664999, 51.84019489438,
    51.8402074312826, 51.8402181772047, 51.8402271321438, 51.8402342960977,
    51.8402396690646, 51.8402432510432, 51.8402450420327, 51.8402450420327,
    51.8402432510432, 51.8402396690646, 51.8402342960977, 51.8402271321438,
    51.8402181772047, 51.8402074312826, 51.84019489438, 51.8401805664999,
    51.8401644476457, 51.8401465378214, 51.8401268370313, 51.8401053452801,
    51.840082062573, 51.8400569889156,
  51.8490481256035, 51.8490732073102, 51.8490964974917, 51.8491179961424,
    51.849137703257, 51.8491556188309, 51.8491717428596, 51.8491860753394,
    51.8491986162667, 51.8492093656387, 51.8492183234525, 51.8492254897062,
    51.849230864398, 51.8492344475266, 51.8492362390911, 51.8492362390911,
    51.8492344475266, 51.849230864398, 51.8492254897062, 51.8492183234525,
    51.8492093656387, 51.8491986162667, 51.8491860753394, 51.8491717428596,
    51.8491556188309, 51.849137703257, 51.8491179961424, 51.8490964974917,
    51.8490732073102, 51.8490481256035,
  51.858039248445, 51.8580643382043, 51.8580876358632, 51.858109141416,
    51.8581288548577, 51.8581467761834, 51.8581629053888, 51.85817724247,
    51.8581897874237, 51.8582005402467, 51.8582095009366, 51.858216669491,
    51.8582220459084, 51.8582256301873, 51.858227422327, 51.858227422327,
    51.8582256301873, 51.8582220459084, 51.858216669491, 51.8582095009366,
    51.8582005402467, 51.8581897874237, 51.85817724247, 51.8581629053888,
    51.8581467761834, 51.8581288548577, 51.858109141416, 51.8580876358632,
    51.8580643382043, 51.858039248445,
  51.8670303574412, 51.8670554552562, 51.8670787603954, 51.8671002728532,
    51.8671199926244, 51.8671379197042, 51.8671540540884, 51.867168395773,
    51.8671809447546, 51.8671917010301, 51.867200664597, 51.8672078354531,
    51.8672132135967, 51.8672167990265, 51.8672185917416, 51.8672185917416,
    51.8672167990265, 51.8672132135967, 51.8672078354531, 51.867200664597,
    51.8671917010301, 51.8671809447546, 51.867168395773, 51.8671540540884,
    51.8671379197042, 51.8671199926244, 51.8671002728532, 51.8670787603954,
    51.8670554552562, 51.8670303574412,
  51.8760214525932, 51.8760465584671, 51.8760698710896, 51.8760913904551,
    51.8761111165583, 51.8761290493946, 51.8761451889595, 51.8761595352493,
    51.8761720882604, 51.8761828479898, 51.8761918144349, 51.8761989875936,
    51.8762043674642, 51.8762079540452, 51.876209747336, 51.876209747336,
    51.8762079540452, 51.8762043674642, 51.8761989875936, 51.8761918144349,
    51.8761828479898, 51.8761720882604, 51.8761595352493, 51.8761451889595,
    51.8761290493946, 51.8761111165583, 51.8760913904551, 51.8760698710896,
    51.8760465584671, 51.8760214525932,
  51.885012533902, 51.8850376478381, 51.8850609679469, 51.8850824942228,
    51.8851022266606, 51.8851201652555, 51.8851363100033, 51.8851506609,
    51.8851632179422, 51.8851739811269, 51.8851829504514, 51.8851901259136,
    51.8851955075118, 51.8851990952446, 51.8852008891112, 51.8852008891112,
    51.8851990952446, 51.8851955075118, 51.8851901259136, 51.8851829504514,
    51.8851739811269, 51.8851632179422, 51.8851506609, 51.8851363100033,
    51.8851201652555, 51.8851022266606, 51.8850824942228, 51.8850609679469,
    51.8850376478381, 51.885012533902,
  51.8940036013687, 51.8940287233701, 51.8940520509682, 51.8940735841573,
    51.8940933229322, 51.8941112672881, 51.8941274172208, 51.8941417727264,
    51.8941543338013, 51.8941651004426, 51.8941740726476, 51.8941812504142,
    51.8941866337407, 51.8941902226257, 51.8941920170684, 51.8941920170684,
    51.8941902226257, 51.8941866337407, 51.8941812504142, 51.8941740726476,
    51.8941651004426, 51.8941543338013, 51.8941417727264, 51.8941274172208,
    51.8941112672881, 51.8940933229322, 51.8940735841573, 51.8940520509682,
    51.8940287233701, 51.8940036013687,
  51.9029946549945, 51.9030197850644, 51.9030431201547, 51.9030646602597,
    51.9030844053742, 51.9031023554935, 51.9031185106131, 51.9031328707293,
    51.9031454358386, 51.9031562059378, 51.9031651810245, 51.9031723610964,
    51.9031777461519, 51.9031813361896, 51.9031831312087, 51.9031831312087,
    51.9031813361896, 51.9031777461519, 51.9031723610964, 51.9031651810245,
    51.9031562059378, 51.9031454358386, 51.9031328707293, 51.9031185106131,
    51.9031023554935, 51.9030844053742, 51.9030646602597, 51.9030431201547,
    51.9030197850644, 51.9029946549945,
  51.9119856947802, 51.912010832922, 51.9120341755075, 51.9120557225312,
    51.9120754739878, 51.9120934298726, 51.9121095901813, 51.91212395491,
    51.9121365240551, 51.9121472976138, 51.9121562755832, 51.9121634579614,
    51.9121688447466, 51.9121724359374, 51.9121742315331, 51.9121742315331,
    51.9121724359374, 51.9121688447466, 51.9121634579614, 51.9121562755832,
    51.9121472976138, 51.9121365240551, 51.91212395491, 51.9121095901813,
    51.9120934298726, 51.9120754739878, 51.9120557225312, 51.9120341755075,
    51.912010832922, 51.9119856947802,
  51.9209767207272, 51.9210018669439, 51.9210252170276, 51.9210467709727,
    51.921066528774, 51.9210844904267, 51.9211006559265, 51.9211150252694,
    51.9211275984521, 51.9211383754715, 51.9211473563249, 51.9211545410103,
    51.9211599295258, 51.9211635218702, 51.9211653180427, 51.9211653180427,
    51.9211635218702, 51.9211599295258, 51.9211545410103, 51.9211473563249,
    51.9211383754715, 51.9211275984521, 51.9211150252694, 51.9211006559265,
    51.9210844904267, 51.921066528774, 51.9210467709727, 51.9210252170276,
    51.9210018669439, 51.9209767207272,
  51.9299677328363, 51.9299928871312, 51.9300162447161, 51.9300378055854,
    51.9300575697338, 51.9300755371567, 51.9300917078497, 51.9301060818088,
    51.9301186590306, 51.9301294395121, 51.9301384232507, 51.9301456102441,
    51.9301510004907, 51.9301545939892, 51.9301563907386, 51.9301563907386,
    51.9301545939892, 51.9301510004907, 51.9301456102441, 51.9301384232507,
    51.9301294395121, 51.9301186590306, 51.9301060818088, 51.9300917078497,
    51.9300755371567, 51.9300575697338, 51.9300378055854, 51.9300162447161,
    51.9299928871312, 51.9299677328363,
  51.9389587311088, 51.9389838934851, 51.9390072585741, 51.9390288263703,
    51.9390485968685, 51.9390665700639, 51.939082745952, 51.9390971245292,
    51.9391097057917, 51.9391204897367, 51.9391294763615, 51.939136665664,
    51.9391420576423, 51.9391456522953, 51.939147449622, 51.939147449622,
    51.9391456522953, 51.9391420576423, 51.939136665664, 51.9391294763615,
    51.9391204897367, 51.9391097057917, 51.9390971245292, 51.939082745952,
    51.9390665700639, 51.9390485968685, 51.9390288263703, 51.9390072585741,
    51.9389838934851, 51.9389587311088,
  51.9479497155456, 51.9479748860065, 51.9479982586027, 51.9480198333287,
    51.9480396101791, 51.9480575891492, 51.9480737702347, 51.9480881534316,
    51.9481007387365, 51.9481115261464, 51.9481205156586, 51.948127707271,
    51.9481331009818, 51.9481366967897, 51.9481384946939, 51.9481384946939,
    51.9481366967897, 51.9481331009818, 51.948127707271, 51.9481205156586,
    51.9481115261464, 51.9481007387365, 51.9480881534316, 51.9480737702347,
    51.9480575891492, 51.9480396101791, 51.9480198333287, 51.9479982586027,
    51.9479748860065, 51.9479497155456,
  51.956940686148, 51.9569658646967, 51.956989244803, 51.9570108264614,
    51.9570306096666, 51.9570485944138, 51.9570647806986, 51.9570791685172,
    51.9570917578661, 51.9571025487423, 51.957111541143, 51.9571187350662,
    51.9571241305102, 51.9571277274735, 51.9571295259554, 51.9571295259554,
    51.9571277274735, 51.9571241305102, 51.9571187350662, 51.957111541143,
    51.9571025487423, 51.9570917578661, 51.9570791685172, 51.9570647806986,
    51.9570485944138, 51.9570306096666, 51.9570108264614, 51.956989244803,
    51.9569658646967, 51.956940686148,
  51.9659316429168, 51.9659568295566, 51.9659802171761, 51.9660018057697,
    51.9660215953322, 51.9660395858587, 51.966055777345, 51.9660701697871,
    51.9660827631816, 51.9660935575254, 51.9661025528158, 51.9661097490508,
    51.9661151462286, 51.9661187443478, 51.9661205434076, 51.9661205434076,
    51.9661187443478, 51.9661151462286, 51.9661097490508, 51.9661025528158,
    51.9660935575254, 51.9660827631816, 51.9660701697871, 51.966055777345,
    51.9660395858587, 51.9660215953322, 51.9660018057697, 51.9659802171761,
    51.9659568295566, 51.9659316429168,
  51.9749225858533, 51.9749477805874, 51.974971175723, 51.9749927712546,
    51.9750125671769, 51.9750305634851, 51.975046760175, 51.9750611572424,
    51.9750737546841, 51.9750845524969, 51.9750935506782, 51.9751007492259,
    51.9751061481381, 51.9751097474137, 51.9751115470517, 51.9751115470517,
    51.9751097474137, 51.9751061481381, 51.9751007492259, 51.9750935506782,
    51.9750845524969, 51.9750737546841, 51.9750611572424, 51.975046760175,
    51.9750305634851, 51.9750125671769, 51.9749927712546, 51.974971175723,
    51.9749477805874, 51.9749225858533,
  51.9839135149585, 51.9839387177901, 51.9839621204449, 51.9839837229172,
    51.9840035252019, 51.9840215272941, 51.9840377291895, 51.9840521308842,
    51.9840647323746, 51.9840755336578, 51.9840845347312, 51.9840917355924,
    51.9840971362399, 51.9841007366723, 51.9841025368887, 51.9841025368887,
    51.9841007366723, 51.9840971362399, 51.9840917355924, 51.9840845347312,
    51.9840755336578, 51.9840647323746, 51.9840521308842, 51.9840377291895,
    51.9840215272941, 51.9840035252019, 51.9839837229172, 51.9839621204449,
    51.9839387177901, 51.9839135149585,
  51.9929044302336, 51.9929296411659, 51.9929530513428, 51.9929746607586,
    51.9929944694082, 51.9930124772867, 51.9930286843898, 51.9930430907135,
    51.9930556962544, 51.9930665010094, 51.9930755049759, 51.9930827081517,
    51.9930881105351, 51.9930917121247, 51.9930935129197, 51.9930935129197,
    51.9930917121247, 51.9930881105351, 51.9930827081517, 51.9930755049759,
    51.9930665010094, 51.9930556962544, 51.9930430907135, 51.9930286843898,
    51.9930124772867, 51.9929944694082, 51.9929746607586, 51.9929530513428,
    51.9929296411659, 51.9929044302336,
  52.0018953316795, 52.0019205507157, 52.0019439684178, 52.0019655847799,
    52.001985399797, 52.0020034134641, 52.0020196257769, 52.0020340367315,
    52.0020466463244, 52.0020574545526, 52.0020664614134, 52.0020736669047,
    52.0020790710246, 52.002082673772, 52.0020844751459, 52.0020844751459,
    52.002082673772, 52.0020790710246, 52.0020736669047, 52.0020664614134,
    52.0020574545526, 52.0020466463244, 52.0020340367315, 52.0020196257769,
    52.0020034134641, 52.001985399797, 52.0019655847799, 52.0019439684178,
    52.0019205507157, 52.0018953316795,
  52.0108862192974, 52.0109114464409, 52.010934871671, 52.0109564949823,
    52.0109763163693, 52.0109943358273, 52.011010553352, 52.0110249689393,
    52.0110375825859, 52.0110483942886, 52.0110574040449, 52.0110646118525,
    52.0110700177098, 52.0110736216153, 52.0110754235684, 52.0110754235684,
    52.0110736216153, 52.0110700177098, 52.0110646118525, 52.0110574040449,
    52.0110483942886, 52.0110375825859, 52.0110249689393, 52.011010553352,
    52.0109943358273, 52.0109763163693, 52.0109564949823, 52.010934871671,
    52.0109114464409, 52.0108862192974,
  52.0198770930883, 52.0199023283423, 52.0199257611036, 52.0199473913667,
    52.0199672191262, 52.0199852443775, 52.020001467116, 52.020015887338,
    52.0200285050398, 52.0200393202185, 52.0200483328714, 52.0200555429964,
    52.0200609505916, 52.0200645556558, 52.0200663581882, 52.0200663581882,
    52.0200645556558, 52.0200609505916, 52.0200555429964, 52.0200483328714,
    52.0200393202185, 52.0200285050398, 52.020015887338, 52.020001467116,
    52.0199852443775, 52.0199672191262, 52.0199473913667, 52.0199257611036,
    52.0199023283423, 52.0198770930883,
  52.0288679530535, 52.0288931964211, 52.0289166367166, 52.0289382739343,
    52.0289581080689, 52.0289761391157, 52.0289923670703, 52.0290067919287,
    52.0290194136874, 52.0290302323434, 52.0290392478941, 52.0290464603373,
    52.0290518696712, 52.0290554758945, 52.0290572790064, 52.0290572790064,
    52.0290554758945, 52.0290518696712, 52.0290464603373, 52.0290392478941,
    52.0290302323434, 52.0290194136874, 52.0290067919287, 52.0289923670703,
    52.0289761391157, 52.0289581080689, 52.0289382739343, 52.0289166367166,
    52.0288931964211, 52.0288679530535,
  52.0378587991939, 52.0378840506785, 52.0379074985112, 52.0379291426862,
    52.0379489831985, 52.0379670200431, 52.0379832532157, 52.0379976827124,
    52.0380103085297, 52.0380211306644, 52.0380301491141, 52.0380373638764,
    52.0380427749497, 52.0380463823326, 52.0380481860243, 52.0380481860243,
    52.0380463823326, 52.0380427749497, 52.0380373638764, 52.0380301491141,
    52.0380211306644, 52.0380103085297, 52.0379976827124, 52.0379832532157,
    52.0379670200431, 52.0379489831985, 52.0379291426862, 52.0379074985112,
    52.0378840506785, 52.0378587991939,
  52.0468496315107, 52.0468748911155, 52.0468983464883, 52.0469199976236,
    52.046939844516, 52.0469578871608, 52.0469741255536, 52.0469885596904,
    52.0470011895678, 52.0470120151827, 52.0470210365324, 52.0470282536148,
    52.0470336664282, 52.0470372749711, 52.0470390792428, 52.0470390792428,
    52.0470372749711, 52.0470336664282, 52.0470282536148, 52.0470210365324,
    52.0470120151827, 52.0470011895678, 52.0469885596904, 52.0469741255536,
    52.0469578871608, 52.046939844516, 52.0469199976236, 52.0468983464883,
    52.0468748911155, 52.0468496315107 ;

 lon =
  4.26478564087425, 4.27928308824974, 4.29378055590363, 4.30827804233386,
    4.32277554603837, 4.33727306551509, 4.35177059926194, 4.36626814577682,
    4.38076570355763, 4.39526327110226, 4.4097608469086, 4.42425842947452,
    4.4387560172979, 4.4532536088766, 4.46775120270851, 4.48224879729149,
    4.49674639112339, 4.5112439827021, 4.52574157052548, 4.5402391530914,
    4.55473672889774, 4.56923429644237, 4.58373185422318, 4.59822940073806,
    4.61272693448491, 4.62722445396163, 4.64172195766614, 4.65621944409637,
    4.67071691175026, 4.68521435912575,
  4.2647438379467, 4.27924416821736, 4.29374451878042, 4.3082448881328,
    4.32274527477138, 4.33724567719307, 4.35174609389473, 4.36624652337324,
    4.38074696412547, 4.39524741464825, 4.40974787343844, 4.42424833899289,
    4.43874880980843, 4.45324928438189, 4.4677497612101, 4.4822502387899,
    4.49675071561811, 4.51125119019157, 4.52575166100711, 4.54025212656156,
    4.55475258535175, 4.56925303587454, 4.58375347662676, 4.59825390610527,
    4.61275432280693, 4.62725472522862, 4.6417551118672, 4.65625548121958,
    4.67075583178264, 4.6852561620533,
  4.26470201322367, 4.27920522789258, 4.29370846286791, 4.30821171664552,
    4.32271498772129, 4.33721827459106, 4.35172157575067, 4.36622488969595,
    4.38072821492273, 4.39523154992682, 4.40973489320404, 4.42423824325017,
    4.43874159856103, 4.45324495763241, 4.4677483189601, 4.4822516810399,
    4.49675504236759, 4.51125840143897, 4.52576175674983, 4.54026510679596,
    4.55476845007318, 4.56927178507727, 4.58377511030405, 4.59827842424933,
    4.61278172540894, 4.62728501227871, 4.64178828335448, 4.65629153713209,
    4.67079477210742, 4.68529798677633,
  4.26466016669011, 4.27916626726138, 4.2936723881531, 4.3081785278601,
    4.3226846848772, 4.33719085769921, 4.35169704482094, 4.36620324473717,
    4.38070945594269, 4.39521567693228, 4.40972190620071, 4.42422814224273,
    4.43873438355312, 4.45324062862662, 4.467746875958, 4.482253124042,
    4.49675937137338, 4.51126561644688, 4.52577185775727, 4.54027809379929,
    4.55478432306772, 4.56929054405731, 4.58379675526283, 4.59830295517907,
    4.61280914230079, 4.6273153151228, 4.6418214721399, 4.6563276118469,
    4.67083373273862, 4.68533983330989,
  4.26461829833095, 4.27912728630974, 4.29363629462301, 4.30814532176457,
    4.32265436622819, 4.33716342650764, 4.35167250109669, 4.36618158848909,
    4.38069068717858, 4.3951997956589, 4.40970891242377, 4.42421803596693,
    4.43872716478209, 4.45323629736297, 4.46774543220327, 4.48225456779673,
    4.49676370263703, 4.51127283521791, 4.52578196403307, 4.54029108757623,
    4.5548002043411, 4.56930931282142, 4.58381841151091, 4.59832749890331,
    4.61283657349236, 4.62734563377181, 4.64185467823543, 4.65636370537699,
    4.67087271369026, 4.68538170166905,
  4.26457640813111, 4.27908828502361, 4.29360018226464, 4.30811209834697,
    4.32262403176334, 4.33713598100647, 4.3516479445691, 4.36615992094392,
    4.38067190862364, 4.39518390610096, 4.40969591186856, 4.42420792441913,
    4.43871994224534, 4.45323196383988, 4.4677439876954, 4.4822560123046,
    4.49676803616012, 4.51128005775466, 4.52579207558087, 4.54030408813144,
    4.55481609389904, 4.56932809137636, 4.58384007905608, 4.5983520554309,
    4.61286401899353, 4.62737596823666, 4.64188790165303, 4.65639981773536,
    4.67091171497639, 4.68542359186889,
  4.2645344960755, 4.27904926338893, 4.29356405106497, 4.30807885759534,
    4.32259368147172, 4.33710852118582, 4.35162337522931, 4.36613824209385,
    4.38065312027111, 4.39516800825273, 4.40968290453038, 4.42419780759568,
    4.43871271594027, 4.45322762805579, 4.46774254243387, 4.48225745756613,
    4.49677237194421, 4.51128728405973, 4.52580219240432, 4.54031709546962,
    4.55483199174727, 4.56934687972889, 4.58386175790615, 4.59837662477069,
    4.61289147881418, 4.62740631852828, 4.64192114240466, 4.65643594893503,
    4.67095073661107, 4.6854655039245,
  4.264492562149, 4.27901022139164, 4.29352790101098, 4.30804559949768,
    4.3225633153424, 4.33708104703578, 4.35159879306845, 4.36611655193106,
    4.3806343221142, 4.39515210210849, 4.40966989040454, 4.42418768549294,
    4.43870548586428, 4.45322329000915, 4.46774109641815, 4.48225890358185,
    4.49677670999085, 4.51129451413572, 4.52581231450707, 4.54033010959546,
    4.55484789789151, 4.5693656778858, 4.58388344806894, 4.59840120693155,
    4.61291895296422, 4.6274366846576, 4.64195440050232, 4.65647209898902,
    4.67098977860836, 4.685507437851,
  4.26445060633649, 4.27897115901766, 4.29349173208962, 4.308012324042,
    4.3225329333644, 4.33705355854643, 4.35157419807768, 4.36609485044772,
    4.38061551414614, 4.3951361876625, 4.40965686948635, 4.42417755810725,
    4.43869825201474, 4.45321894969839, 4.46773964964772, 4.48226035035228,
    4.49678105030161, 4.51130174798525, 4.52582244189275, 4.54034313051365,
    4.5548638123375, 4.56938448585386, 4.58390514955228, 4.59842580192232,
    4.61294644145357, 4.6274670666356, 4.641987675958, 4.65650826791038,
    4.67102884098234, 4.68554939366351,
  4.26440862862282, 4.27893207625289, 4.29345554428785, 4.30797903121629,
    4.32250253552678, 4.33702605570787, 4.3515495902481, 4.36607313763602,
    4.38059669636015, 4.395120264909, 4.4096438417711, 4.42416742543496,
    4.43869101438907, 4.45321460712194, 4.46773820212206, 4.48226179787794,
    4.49678539287806, 4.51130898561093, 4.52583257456504, 4.5403561582289,
    4.554879735091, 4.56940330363985, 4.58392686236398, 4.5984504097519,
    4.61297394429213, 4.62749746447322, 4.64202096878371, 4.65654445571215,
    4.67106792374711, 4.68559137137718,
  4.26436662899285, 4.27889297308321, 4.2934193375926, 4.30794572100854,
    4.32247212181856, 4.33699853851016, 4.35152496957084, 4.3660514134881,
    4.38057786874942, 4.39510433384226, 4.40963080725411, 4.42415728747241,
    4.43868377298464, 4.45321026227823, 4.46773675384065, 4.48226324615935,
    4.49678973772177, 4.51131622701536, 4.52584271252759, 4.54036919274589,
    4.55489566615774, 4.56942213125058, 4.5839485865119, 4.59847503042916,
    4.61300146148984, 4.62752787818144, 4.64205427899146, 4.6565806624074,
    4.67110702691679, 4.68563337100715,
  4.2643246074314, 4.27885384949452, 4.29338311199079, 4.30791239340671,
    4.32244169222875, 4.33697100694336, 4.35150033603701, 4.36602967799613,
    4.38055903130716, 4.39508839445653, 4.40961776593065, 4.42414714421595,
    4.43867652779883, 4.4532059151657, 4.46773530480297, 4.48226469519703,
    4.4967940848343, 4.51132347220117, 4.52585285578405, 4.54038223406935,
    4.55491160554347, 4.56944096869284, 4.58397032200387, 4.59849966396299,
    4.61302899305664, 4.62755830777125, 4.64208760659329, 4.65661688800921,
    4.67114615050548, 4.6856753925686,
  4.2642825639233, 4.27881470547267, 4.29334686746934, 4.30787904839877,
    4.32241124674635, 4.33694346099753, 4.3514756896377, 4.36600793115224,
    4.38054018402656, 4.39507244674603, 4.40960471779602, 4.4241369956619,
    4.43866927882903, 4.45320156578277, 4.46773385500848, 4.48226614499152,
    4.49679843421723, 4.51133072117097, 4.5258630043381, 4.54039528220398,
    4.55492755325397, 4.56945981597344, 4.58399206884776, 4.5985243103623,
    4.61305653900247, 4.62758875325364, 4.64212095160123, 4.65665313253066,
    4.67118529452733, 4.6857174360767,
  4.26424049845334, 4.27877554100351, 4.29331060401515, 4.30784568597265,
    4.32238078536038, 4.33691590066271, 4.351451030364, 4.36598617294859,
    4.38052132690082, 4.39505649070501, 4.4095916628455, 4.4241268418066,
    4.43866202607262, 4.45319721412788, 4.46773240445668, 4.48226759554332,
    4.49680278587212, 4.51133797392738, 4.5258731581934, 4.5404083371545,
    4.55494350929499, 4.56947867309918, 4.58401382705141, 4.598548969636,
    4.61308409933729, 4.62761921463962, 4.64215431402735, 4.65668939598485,
    4.67122445899649, 4.68575950154667,
  4.26419841100631, 4.27873635607288, 4.29327432161509, 4.30781230611629,
    4.3223503080598, 4.33688832592893, 4.351426358207, 4.36596440337729,
    4.3805024599231, 4.3950405263277, 4.40957860107437, 4.42411668264638,
    4.43865476952698, 4.45319286019944, 4.46773095314702, 4.48226904685298,
    4.49680713980056, 4.51134523047302, 4.52588331735362, 4.54042139892563,
    4.5549594736723, 4.5694975400769, 4.58403559662271, 4.598573641793,
    4.61311167407107, 4.6276496919402, 4.64218769388371, 4.65672567838491,
    4.67126364392712, 4.68580158899369,
  4.26415630156699, 4.2786971506666, 4.29323802025605, 4.30777890881762,
    4.32231981483359, 4.33686073678622, 4.35140167315777, 4.36594262243048,
    4.38048358308659, 4.39502455360832, 4.4095655324779, 4.42410651817755,
    4.43864750918948, 4.45318850399589, 4.467729501079, 4.482270498921,
    4.49681149600411, 4.51135249081052, 4.52589348182245, 4.5404344675221,
    4.55497544639168, 4.56951641691341, 4.58405737756952, 4.59859832684223,
    4.61313926321378, 4.62768018516641, 4.64222109118238, 4.65676197974395,
    4.6713028493334, 4.68584369843301,
  4.26411417012013, 4.27865792477049, 4.29320169992489, 4.30774549406455,
    4.32228930567072, 4.33683313322459, 4.35137697520738, 4.36592083010027,
    4.38046469638445, 4.39500857254109, 4.40955245705137, 4.42409634839645,
    4.43864024505749, 4.45318414551565, 4.46772804825207, 4.48227195174793,
    4.49681585448435, 4.51135975494251, 4.52590365160355, 4.54044754294863,
    4.55499142745891, 4.56953530361555, 4.58407916989973, 4.59862302479262,
    4.61316686677541, 4.62771069432928, 4.64225450593545, 4.65679830007511,
    4.67134207522951, 4.68588582987987,
  4.26407201665049, 4.27861867837034, 4.29316536060845, 4.30771206184499,
    4.32225878056013, 4.33680551523405, 4.35135226434688, 4.36589902637877,
    4.38044579980984, 4.39499258312022, 4.40953937479004, 4.42408617329939,
    4.43863297712838, 4.45317978475713, 4.46772659466573, 4.48227340533427,
    4.49682021524287, 4.51136702287162, 4.52591382670061, 4.54046062520996,
    4.55500741687978, 4.56955420019016, 4.58410097362123, 4.59864773565312,
    4.61319448476595, 4.62774121943987, 4.64228793815501, 4.65683463939155,
    4.67138132162966, 4.68592798334951,
  4.26402984114279, 4.27857941145194, 4.29312900229357, 4.30767861214681,
    4.32222823949078, 4.33677788280459, 4.35132754056732, 4.36587721125808,
    4.38042689335592, 4.39497658533993, 4.40952628568916, 4.42407599288267,
    4.43862570539953, 4.45317542171876, 4.46772514031943, 4.48227485968057,
    4.49682457828124, 4.51137429460047, 4.52592400711733, 4.54047371431084,
    4.55502341466007, 4.56957310664408, 4.58412278874192, 4.59867245943268,
    4.61322211719541, 4.62777176050922, 4.64232138785319, 4.65687099770643,
    4.67142058854806, 4.68597015885721,
  4.26398764358175, 4.27854012400105, 4.29309262496708, 4.3076451449579,
    4.32219768245159, 4.3367502359262, 4.35130280385975, 4.36585538473029,
    4.38040797701584, 4.39496057919441, 4.409513189744, 4.42406580714263,
    4.43861842986828, 4.45317105639896, 4.46772368521265, 4.48227631478735,
    4.49682894360104, 4.51138157013172, 4.52593419285737, 4.540486810256,
    4.55503942080559, 4.56959202298416, 4.5841446152697, 4.59869719614025,
    4.6132497640738, 4.62780231754841, 4.6423548550421, 4.65690737503292,
    4.67145987599895, 4.68601235641825,
  4.26394542395207, 4.27850081600343, 4.29305622861578, 4.30761166026613,
    4.32216710943149, 4.33672257458885, 4.3512780542152, 4.3658335467875,
    4.38038905078274, 4.39494456467786, 4.40950008694981, 4.42405561607555,
    4.43861115053202, 4.45316668879614, 4.46772222934487, 4.48227777065513,
    4.49683331120386, 4.51138884946798, 4.52594438392445, 4.54049991305019,
    4.55505543532214, 4.56961094921726, 4.5841664532125, 4.5987219457848,
    4.61327742541115, 4.62783289056851, 4.64238833973387, 4.65694377138422,
    4.67149918399657, 4.68605457604793,
  4.26390318223843, 4.27846148744483, 4.29301981322648, 4.30757815805935,
    4.32213652041938, 4.33669489878251, 4.35125329162468, 4.36581169742179,
    4.38037011464975, 4.39492854178447, 4.40948697730184, 4.42404541967775,
    4.43860386738809, 4.45316231890873, 4.46772077271556, 4.48227922728444,
    4.49683768109127, 4.51139613261191, 4.52595458032225, 4.54051302269816,
    4.55507145821553, 4.56962988535025, 4.58418830257821, 4.59874670837532,
    4.61330510121749, 4.62786347958062, 4.64242184194065, 4.65698018677352,
    4.67153851255517, 4.68609681776157,
  4.26386091842551, 4.27842213831097, 4.29298337878596, 4.3075446383254,
    4.32210591540417, 4.33666720849715, 4.35122851607921, 4.36578983662521,
    4.38035116861001, 4.39491251050843, 4.40947386079533, 4.42403521794553,
    4.43859658043385, 4.45315794673513, 4.46771931532418, 4.48228068467582,
    4.49684205326487, 4.51140341956615, 4.52596478205447, 4.54052613920467,
    4.55508748949157, 4.56964883139, 4.58421016337479, 4.59877148392079,
    4.61333279150285, 4.62789408459583, 4.6424553616746, 4.65701662121404,
    4.67157786168903, 4.68613908157449,
  4.26381863249797, 4.27838276858757, 4.292946925281, 4.30751110105212,
    4.32207529437474, 4.3366395037227, 4.3512037275698, 4.36576796438985,
    4.38033221265662, 4.39489647084392, 4.40946073742551, 4.42402501087517,
    4.43858928966667, 4.45315357227376, 4.46771785717021, 4.48228214282979,
    4.49684642772624, 4.51141071033333, 4.52597498912483, 4.54053926257449,
    4.55510352915608, 4.56966778734338, 4.58423203561015, 4.5987962724302,
    4.6133604962773, 4.62792470562526, 4.64248889894788, 4.657053074719,
    4.67161723141243, 4.68618136750203,
  4.26377632444045, 4.27834337826033, 4.29291045269836, 4.30747754622732,
    4.32204465731998, 4.33661178444911, 4.35117892608745, 4.36574608070775,
    4.38031324678272, 4.39488042278511, 4.40944760718763, 4.42401479846298,
    4.43858199508388, 4.45314919552303, 4.46771639825312, 4.48228360174687,
    4.49685080447697, 4.51141800491612, 4.52598520153702, 4.54055239281237,
    4.55511957721489, 4.56968675321728, 4.58425391929226, 4.59882107391255,
    4.61338821555089, 4.62795534268002, 4.64252245377268, 4.65708954730164,
    4.67165662173967, 4.68622367555955,
  4.26373399423758, 4.27830396731494, 4.29287396102478, 4.30744397383882,
    4.32201400422876, 4.3365840506663, 4.35115411162314, 4.36572418557096,
    4.38029427098141, 4.39486436632618, 4.4094344700769, 4.42400458070524,
    4.43857469668284, 4.45314481648134, 4.46771493857239, 4.48228506142761,
    4.49685518351866, 4.51142530331716, 4.52599541929476, 4.5405655299231,
    4.55513563367382, 4.56970572901859, 4.58427581442904, 4.59884588837686,
    4.6134159493337, 4.62798599577124, 4.64255602616118, 4.65712603897522,
    4.67169603268505, 4.68626600576242,
  4.26369164187397, 4.27826453573708, 4.29283745024701, 4.30741038387441,
    4.32198333508992, 4.3365563023642, 4.35112928416786, 4.36570227897152,
    4.3802752852458, 4.39484830146128, 4.40942132608857, 4.42399435759825,
    4.4385673944609, 4.45314043514712, 4.46771347812747, 4.48228652187253,
    4.49685956485288, 4.5114326055391, 4.52600564240175, 4.54057867391143,
    4.55515169853872, 4.5697247147542, 4.58429772102848, 4.59887071583214,
    4.6134436976358, 4.62801666491008, 4.64258961612559, 4.65716254975299,
    4.67173546426292, 4.68630835812603,
  4.26364926733422, 4.27822508351241, 4.29280092035176, 4.30737677632187,
    4.32195264989233, 4.33652853953271, 4.35110444371258, 4.36568036090148,
    4.38025628956897, 4.39483222818458, 4.40940817521783, 4.42398412913827,
    4.43856008841541, 4.45313605151876, 4.46771201691784, 4.48228798308216,
    4.49686394848124, 4.51143991158459, 4.52601587086173, 4.54059182478217,
    4.55516777181542, 4.56974371043103, 4.58431963909852, 4.59889555628742,
    4.61347146046729, 4.62804735010767, 4.64262322367813, 4.65719907964824,
    4.67177491648759, 4.68635073266578,
  4.26360687060292, 4.27818561062657, 4.29276437132575, 4.30734315116899,
    4.32192194862482, 4.33650076216174, 4.35107959024825, 4.36565843135285,
    4.38023728394402, 4.39481614649022, 4.40939501745992, 4.4239738953216,
    4.43855277854369, 4.45313166559467, 4.46771055494296, 4.48228944505704,
    4.49686833440533, 4.51144722145631, 4.5260261046784, 4.54060498254008,
    4.55518385350978, 4.56976271605598, 4.58434156864715, 4.59892040975175,
    4.61349923783826, 4.62807805137518, 4.64265684883101, 4.65723562867425,
    4.67181438937343, 4.68639312939708,
  4.26356445166463, 4.2781461170652, 4.29272780315567, 4.30730950840352,
    4.3218912312762, 4.33647297024117, 4.35105472376584, 4.36563649031766,
    4.38021826836403, 4.39480005637236, 4.40938185281005, 4.4239636561445,
    4.4385454648431, 4.45312727737325, 4.46770909220231, 4.48229090779769,
    4.49687272262675, 4.5114545351569, 4.5260363438555, 4.54061814718995,
    4.55519994362764, 4.56978173163597, 4.58436350968234, 4.59894527623416,
    4.61352702975883, 4.6281087687238, 4.64269049159648, 4.65727219684433,
    4.6718538829348, 4.68643554833537 ;

 rlat = 51.914378775434, 51.9089235868341, 51.9280541060936,
    51.9221924255006, 51.8675636655372, 51.9329093410371, 51.9374470181688,
    51.8702273745715, 51.9569447692371 ;

 rlon = 4.48023556929616, 4.32489363985269, 4.4616468480345,
    4.40183718531446, 4.35517721897712, 4.22860389049183, 4.43333892655883,
    4.58046723703735, 4.43722152827864 ;

 weights = 0.142857142857143, 0.142857142857143, 0.142857142857143,
    0.142857142857143, 0.142857142857143, 0.142857142857143, 0.142857142857143 ;
}
